----------------------------------------------
-- Erzeugt mit Create_Blockram
--   InFilename   = ..\Software\TestDMA\Debug\TestDMA.hex
--   Templatename = template_bsr2_rom.vhd
--   Startadresse = 0x0
--   Endadresse   = 0x37ff
-- (Prof. Bernhard Lang, FH Osnabrueck)
----------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bsr2_rom is
 port(
  CLK_I  : in  std_logic;
  RST_I  : in  std_logic;
  STB_I  : in  std_logic;
  WE_I   : in  std_logic;
  SEL_I  : in  std_logic_vector(3 downto 0);
  ADR_I  : in  std_logic_vector(13 downto 0);
  DAT_I  : in  std_logic_vector(31 downto 0);
  DAT_O  : out std_logic_vector(31 downto 0);
  ACK_O  : out std_logic
  );
end entity;

architecture behavioral of bsr2_rom is
  type memory_t is array (0 to 2 ** (ADR_I'length - 2) - 1) of std_logic_vector(31 downto 0);

  signal read_ack  : std_logic := '0';
  signal write_ack : std_logic;
  signal DAT_O_i   : std_logic_vector(31 downto 0) := (others=>'-');
  signal memory    : memory_t := (
    x"10000013", -- 0x00000000
    x"00000000", -- 0x00000004
    x"00000000", -- 0x00000008
    x"00000000", -- 0x0000000c
    x"10000017", -- 0x00000010
    x"00000000", -- 0x00000014
    x"00000000", -- 0x00000018
    x"00000000", -- 0x0000001c
    x"1000001b", -- 0x00000020
    x"00000000", -- 0x00000024
    x"00000000", -- 0x00000028
    x"00000000", -- 0x0000002c
    x"1000001f", -- 0x00000030
    x"00000000", -- 0x00000034
    x"00000000", -- 0x00000038
    x"00000000", -- 0x0000003c
    x"10000023", -- 0x00000040
    x"00000000", -- 0x00000044
    x"00000000", -- 0x00000048
    x"00000000", -- 0x0000004c
    x"3c1d0001", -- 0x00000050
    x"27bd8000", -- 0x00000054
    x"3c1e0001", -- 0x00000058
    x"27de8000", -- 0x0000005c
    x"3c1c0000", -- 0x00000060
    x"279c4000", -- 0x00000064
    x"41606020", -- 0x00000068
    x"08000493", -- 0x0000006c
    x"27bdffb8", -- 0x00000070
    x"afbf0000", -- 0x00000074
    x"0c00003c", -- 0x00000078
    x"0c000146", -- 0x0000007c
    x"0c00004e", -- 0x00000080
    x"8fbf0000", -- 0x00000084
    x"27bd0048", -- 0x00000088
    x"42000018", -- 0x0000008c
    x"27bdffb8", -- 0x00000090
    x"afbf0000", -- 0x00000094
    x"0c00003c", -- 0x00000098
    x"0c000362", -- 0x0000009c
    x"0c00004e", -- 0x000000a0
    x"8fbf0000", -- 0x000000a4
    x"27bd0048", -- 0x000000a8
    x"42000018", -- 0x000000ac
    x"27bdffb8", -- 0x000000b0
    x"afbf0000", -- 0x000000b4
    x"0c00003c", -- 0x000000b8
    x"0c000158", -- 0x000000bc
    x"0c00004e", -- 0x000000c0
    x"8fbf0000", -- 0x000000c4
    x"27bd0048", -- 0x000000c8
    x"42000018", -- 0x000000cc
    x"27bdffb8", -- 0x000000d0
    x"afbf0000", -- 0x000000d4
    x"0c00003c", -- 0x000000d8
    x"0c000161", -- 0x000000dc
    x"0c00004e", -- 0x000000e0
    x"8fbf0000", -- 0x000000e4
    x"27bd0048", -- 0x000000e8
    x"42000018", -- 0x000000ec
    x"afa10004", -- 0x000000f0
    x"afa20008", -- 0x000000f4
    x"afa3000c", -- 0x000000f8
    x"afa40010", -- 0x000000fc
    x"afa50014", -- 0x00000100
    x"afa60018", -- 0x00000104
    x"afa7001c", -- 0x00000108
    x"afa80020", -- 0x0000010c
    x"afa90024", -- 0x00000110
    x"afaa0028", -- 0x00000114
    x"afab002c", -- 0x00000118
    x"afac0030", -- 0x0000011c
    x"afad0034", -- 0x00000120
    x"afae0038", -- 0x00000124
    x"afaf003c", -- 0x00000128
    x"afb80040", -- 0x0000012c
    x"afb90044", -- 0x00000130
    x"03e00008", -- 0x00000134
    x"8fa10004", -- 0x00000138
    x"8fa20008", -- 0x0000013c
    x"8fa3000c", -- 0x00000140
    x"8fa40010", -- 0x00000144
    x"8fa50014", -- 0x00000148
    x"8fa60018", -- 0x0000014c
    x"8fa7001c", -- 0x00000150
    x"8fa80020", -- 0x00000154
    x"8fa90024", -- 0x00000158
    x"8faa0028", -- 0x0000015c
    x"8fab002c", -- 0x00000160
    x"8fac0030", -- 0x00000164
    x"8fad0034", -- 0x00000168
    x"8fae0038", -- 0x0000016c
    x"8faf003c", -- 0x00000170
    x"8fb80040", -- 0x00000174
    x"8fb90044", -- 0x00000178
    x"03e00008", -- 0x0000017c
    x"41626020", -- 0x00000180
    x"03e00008", -- 0x00000184
    x"41626000", -- 0x00000188
    x"03e00008", -- 0x0000018c
    x"27bdfff8", -- 0x00000190
    x"afbe0004", -- 0x00000194
    x"03a0f025", -- 0x00000198
    x"afc40008", -- 0x0000019c
    x"afc5000c", -- 0x000001a0
    x"afc60010", -- 0x000001a4
    x"8fc20008", -- 0x000001a8
    x"00000000", -- 0x000001ac
    x"ac400000", -- 0x000001b0
    x"8fc20008", -- 0x000001b4
    x"00000000", -- 0x000001b8
    x"ac400004", -- 0x000001bc
    x"8fc20008", -- 0x000001c0
    x"8fc30010", -- 0x000001c4
    x"00000000", -- 0x000001c8
    x"ac430008", -- 0x000001cc
    x"8fc20008", -- 0x000001d0
    x"8fc3000c", -- 0x000001d4
    x"00000000", -- 0x000001d8
    x"ac43000c", -- 0x000001dc
    x"00000000", -- 0x000001e0
    x"03c0e825", -- 0x000001e4
    x"8fbe0004", -- 0x000001e8
    x"27bd0008", -- 0x000001ec
    x"03e00008", -- 0x000001f0
    x"00000000", -- 0x000001f4
    x"27bdfff0", -- 0x000001f8
    x"afbe000c", -- 0x000001fc
    x"03a0f025", -- 0x00000200
    x"afc40010", -- 0x00000204
    x"afc50014", -- 0x00000208
    x"8fc20010", -- 0x0000020c
    x"00000000", -- 0x00000210
    x"8c430000", -- 0x00000214
    x"8fc20010", -- 0x00000218
    x"00000000", -- 0x0000021c
    x"8c420004", -- 0x00000220
    x"00000000", -- 0x00000224
    x"00621023", -- 0x00000228
    x"2442ffff", -- 0x0000022c
    x"afc20000", -- 0x00000230
    x"8fc20000", -- 0x00000234
    x"00000000", -- 0x00000238
    x"04410008", -- 0x0000023c
    x"00000000", -- 0x00000240
    x"8fc20010", -- 0x00000244
    x"00000000", -- 0x00000248
    x"8c430008", -- 0x0000024c
    x"8fc20000", -- 0x00000250
    x"00000000", -- 0x00000254
    x"00621021", -- 0x00000258
    x"afc20000", -- 0x0000025c
    x"8fc20000", -- 0x00000260
    x"00000000", -- 0x00000264
    x"18400034", -- 0x00000268
    x"00000000", -- 0x0000026c
    x"8fc20010", -- 0x00000270
    x"00000000", -- 0x00000274
    x"8c42000c", -- 0x00000278
    x"8fc30010", -- 0x0000027c
    x"00000000", -- 0x00000280
    x"8c630004", -- 0x00000284
    x"00000000", -- 0x00000288
    x"00431021", -- 0x0000028c
    x"8fc30014", -- 0x00000290
    x"00000000", -- 0x00000294
    x"306300ff", -- 0x00000298
    x"a0430000", -- 0x0000029c
    x"8fc20010", -- 0x000002a0
    x"00000000", -- 0x000002a4
    x"8c420004", -- 0x000002a8
    x"00000000", -- 0x000002ac
    x"24430001", -- 0x000002b0
    x"8fc20010", -- 0x000002b4
    x"00000000", -- 0x000002b8
    x"ac430004", -- 0x000002bc
    x"8fc20010", -- 0x000002c0
    x"00000000", -- 0x000002c4
    x"8c420004", -- 0x000002c8
    x"00000000", -- 0x000002cc
    x"00401825", -- 0x000002d0
    x"8fc20010", -- 0x000002d4
    x"00000000", -- 0x000002d8
    x"8c420008", -- 0x000002dc
    x"00000000", -- 0x000002e0
    x"0062102b", -- 0x000002e4
    x"1440000f", -- 0x000002e8
    x"00000000", -- 0x000002ec
    x"8fc20010", -- 0x000002f0
    x"00000000", -- 0x000002f4
    x"8c420004", -- 0x000002f8
    x"00000000", -- 0x000002fc
    x"00401825", -- 0x00000300
    x"8fc20010", -- 0x00000304
    x"00000000", -- 0x00000308
    x"8c420008", -- 0x0000030c
    x"00000000", -- 0x00000310
    x"00621023", -- 0x00000314
    x"00401825", -- 0x00000318
    x"8fc20010", -- 0x0000031c
    x"00000000", -- 0x00000320
    x"ac430004", -- 0x00000324
    x"8fc20000", -- 0x00000328
    x"00000000", -- 0x0000032c
    x"2442ffff", -- 0x00000330
    x"10000002", -- 0x00000334
    x"00000000", -- 0x00000338
    x"2402ffff", -- 0x0000033c
    x"03c0e825", -- 0x00000340
    x"8fbe000c", -- 0x00000344
    x"27bd0010", -- 0x00000348
    x"03e00008", -- 0x0000034c
    x"00000000", -- 0x00000350
    x"27bdfff0", -- 0x00000354
    x"afbe000c", -- 0x00000358
    x"03a0f025", -- 0x0000035c
    x"afc40010", -- 0x00000360
    x"afc50014", -- 0x00000364
    x"8fc20010", -- 0x00000368
    x"00000000", -- 0x0000036c
    x"8c430004", -- 0x00000370
    x"8fc20010", -- 0x00000374
    x"00000000", -- 0x00000378
    x"8c420000", -- 0x0000037c
    x"00000000", -- 0x00000380
    x"00621023", -- 0x00000384
    x"afc20000", -- 0x00000388
    x"8fc20000", -- 0x0000038c
    x"00000000", -- 0x00000390
    x"04410008", -- 0x00000394
    x"00000000", -- 0x00000398
    x"8fc20010", -- 0x0000039c
    x"00000000", -- 0x000003a0
    x"8c430008", -- 0x000003a4
    x"8fc20000", -- 0x000003a8
    x"00000000", -- 0x000003ac
    x"00621021", -- 0x000003b0
    x"afc20000", -- 0x000003b4
    x"8fc20000", -- 0x000003b8
    x"00000000", -- 0x000003bc
    x"18400034", -- 0x000003c0
    x"00000000", -- 0x000003c4
    x"8fc20010", -- 0x000003c8
    x"00000000", -- 0x000003cc
    x"8c42000c", -- 0x000003d0
    x"8fc30010", -- 0x000003d4
    x"00000000", -- 0x000003d8
    x"8c630000", -- 0x000003dc
    x"00000000", -- 0x000003e0
    x"00431021", -- 0x000003e4
    x"90430000", -- 0x000003e8
    x"8fc20014", -- 0x000003ec
    x"00000000", -- 0x000003f0
    x"a0430000", -- 0x000003f4
    x"8fc20010", -- 0x000003f8
    x"00000000", -- 0x000003fc
    x"8c420000", -- 0x00000400
    x"00000000", -- 0x00000404
    x"24430001", -- 0x00000408
    x"8fc20010", -- 0x0000040c
    x"00000000", -- 0x00000410
    x"ac430000", -- 0x00000414
    x"8fc20010", -- 0x00000418
    x"00000000", -- 0x0000041c
    x"8c420000", -- 0x00000420
    x"00000000", -- 0x00000424
    x"00401825", -- 0x00000428
    x"8fc20010", -- 0x0000042c
    x"00000000", -- 0x00000430
    x"8c420008", -- 0x00000434
    x"00000000", -- 0x00000438
    x"0062102b", -- 0x0000043c
    x"1440000f", -- 0x00000440
    x"00000000", -- 0x00000444
    x"8fc20010", -- 0x00000448
    x"00000000", -- 0x0000044c
    x"8c420000", -- 0x00000450
    x"00000000", -- 0x00000454
    x"00401825", -- 0x00000458
    x"8fc20010", -- 0x0000045c
    x"00000000", -- 0x00000460
    x"8c420008", -- 0x00000464
    x"00000000", -- 0x00000468
    x"00621023", -- 0x0000046c
    x"00401825", -- 0x00000470
    x"8fc20010", -- 0x00000474
    x"00000000", -- 0x00000478
    x"ac430000", -- 0x0000047c
    x"8fc20000", -- 0x00000480
    x"00000000", -- 0x00000484
    x"2442ffff", -- 0x00000488
    x"10000002", -- 0x0000048c
    x"00000000", -- 0x00000490
    x"2402ffff", -- 0x00000494
    x"03c0e825", -- 0x00000498
    x"8fbe000c", -- 0x0000049c
    x"27bd0010", -- 0x000004a0
    x"03e00008", -- 0x000004a4
    x"00000000", -- 0x000004a8
    x"27bdfff8", -- 0x000004ac
    x"afbe0004", -- 0x000004b0
    x"03a0f025", -- 0x000004b4
    x"afc40008", -- 0x000004b8
    x"afc5000c", -- 0x000004bc
    x"8fc20008", -- 0x000004c0
    x"8fc3000c", -- 0x000004c4
    x"00000000", -- 0x000004c8
    x"ac430000", -- 0x000004cc
    x"00000000", -- 0x000004d0
    x"03c0e825", -- 0x000004d4
    x"8fbe0004", -- 0x000004d8
    x"27bd0008", -- 0x000004dc
    x"03e00008", -- 0x000004e0
    x"00000000", -- 0x000004e4
    x"27bdfff8", -- 0x000004e8
    x"afbe0004", -- 0x000004ec
    x"03a0f025", -- 0x000004f0
    x"afc40008", -- 0x000004f4
    x"8fc20008", -- 0x000004f8
    x"00000000", -- 0x000004fc
    x"8c420000", -- 0x00000500
    x"03c0e825", -- 0x00000504
    x"8fbe0004", -- 0x00000508
    x"27bd0008", -- 0x0000050c
    x"03e00008", -- 0x00000510
    x"00000000", -- 0x00000514
    x"27bdfff8", -- 0x00000518
    x"afbe0004", -- 0x0000051c
    x"03a0f025", -- 0x00000520
    x"00000000", -- 0x00000524
    x"03c0e825", -- 0x00000528
    x"8fbe0004", -- 0x0000052c
    x"27bd0008", -- 0x00000530
    x"03e00008", -- 0x00000534
    x"00000000", -- 0x00000538
    x"27bdfff8", -- 0x0000053c
    x"afbe0004", -- 0x00000540
    x"03a0f025", -- 0x00000544
    x"00000000", -- 0x00000548
    x"03c0e825", -- 0x0000054c
    x"8fbe0004", -- 0x00000550
    x"27bd0008", -- 0x00000554
    x"03e00008", -- 0x00000558
    x"00000000", -- 0x0000055c
    x"27bdfff8", -- 0x00000560
    x"afbe0004", -- 0x00000564
    x"03a0f025", -- 0x00000568
    x"00000000", -- 0x0000056c
    x"03c0e825", -- 0x00000570
    x"8fbe0004", -- 0x00000574
    x"27bd0008", -- 0x00000578
    x"03e00008", -- 0x0000057c
    x"00000000", -- 0x00000580
    x"27bdfff8", -- 0x00000584
    x"afbe0004", -- 0x00000588
    x"03a0f025", -- 0x0000058c
    x"00000000", -- 0x00000590
    x"03c0e825", -- 0x00000594
    x"8fbe0004", -- 0x00000598
    x"27bd0008", -- 0x0000059c
    x"03e00008", -- 0x000005a0
    x"00000000", -- 0x000005a4
    x"27bdffe0", -- 0x000005a8
    x"afbf001c", -- 0x000005ac
    x"afbe0018", -- 0x000005b0
    x"03a0f025", -- 0x000005b4
    x"afc40020", -- 0x000005b8
    x"2404000c", -- 0x000005bc
    x"0c00019c", -- 0x000005c0
    x"00000000", -- 0x000005c4
    x"afc20010", -- 0x000005c8
    x"8fc30010", -- 0x000005cc
    x"8fc20020", -- 0x000005d0
    x"00000000", -- 0x000005d4
    x"00621025", -- 0x000005d8
    x"00402825", -- 0x000005dc
    x"2404000c", -- 0x000005e0
    x"0c0001bf", -- 0x000005e4
    x"00000000", -- 0x000005e8
    x"00000000", -- 0x000005ec
    x"03c0e825", -- 0x000005f0
    x"8fbf001c", -- 0x000005f4
    x"8fbe0018", -- 0x000005f8
    x"27bd0020", -- 0x000005fc
    x"03e00008", -- 0x00000600
    x"00000000", -- 0x00000604
    x"27bdffe0", -- 0x00000608
    x"afbf001c", -- 0x0000060c
    x"afbe0018", -- 0x00000610
    x"03a0f025", -- 0x00000614
    x"afc40020", -- 0x00000618
    x"2404000c", -- 0x0000061c
    x"0c00019c", -- 0x00000620
    x"00000000", -- 0x00000624
    x"afc20010", -- 0x00000628
    x"8fc20020", -- 0x0000062c
    x"00000000", -- 0x00000630
    x"00021827", -- 0x00000634
    x"8fc20010", -- 0x00000638
    x"00000000", -- 0x0000063c
    x"00621024", -- 0x00000640
    x"00402825", -- 0x00000644
    x"2404000c", -- 0x00000648
    x"0c0001bf", -- 0x0000064c
    x"00000000", -- 0x00000650
    x"00000000", -- 0x00000654
    x"03c0e825", -- 0x00000658
    x"8fbf001c", -- 0x0000065c
    x"8fbe0018", -- 0x00000660
    x"27bd0020", -- 0x00000664
    x"03e00008", -- 0x00000668
    x"00000000", -- 0x0000066c
    x"27bdfff0", -- 0x00000670
    x"afbe000c", -- 0x00000674
    x"03a0f025", -- 0x00000678
    x"afc40010", -- 0x0000067c
    x"afc00000", -- 0x00000680
    x"8fc20010", -- 0x00000684
    x"2403000d", -- 0x00000688
    x"1043000c", -- 0x0000068c
    x"00000000", -- 0x00000690
    x"2403000e", -- 0x00000694
    x"1043000e", -- 0x00000698
    x"00000000", -- 0x0000069c
    x"2403000c", -- 0x000006a0
    x"1443000f", -- 0x000006a4
    x"00000000", -- 0x000006a8
    x"40026000", -- 0x000006ac
    x"00000000", -- 0x000006b0
    x"afc20000", -- 0x000006b4
    x"1000000a", -- 0x000006b8
    x"00000000", -- 0x000006bc
    x"40026800", -- 0x000006c0
    x"00000000", -- 0x000006c4
    x"afc20000", -- 0x000006c8
    x"10000005", -- 0x000006cc
    x"00000000", -- 0x000006d0
    x"40027000", -- 0x000006d4
    x"00000000", -- 0x000006d8
    x"afc20000", -- 0x000006dc
    x"00000000", -- 0x000006e0
    x"8fc20000", -- 0x000006e4
    x"03c0e825", -- 0x000006e8
    x"8fbe000c", -- 0x000006ec
    x"27bd0010", -- 0x000006f0
    x"03e00008", -- 0x000006f4
    x"00000000", -- 0x000006f8
    x"27bdfff8", -- 0x000006fc
    x"afbe0004", -- 0x00000700
    x"03a0f025", -- 0x00000704
    x"afc40008", -- 0x00000708
    x"afc5000c", -- 0x0000070c
    x"8fc20008", -- 0x00000710
    x"2403000d", -- 0x00000714
    x"1043000e", -- 0x00000718
    x"00000000", -- 0x0000071c
    x"2403000e", -- 0x00000720
    x"10430010", -- 0x00000724
    x"00000000", -- 0x00000728
    x"2403000c", -- 0x0000072c
    x"10430003", -- 0x00000730
    x"00000000", -- 0x00000734
    x"1000000f", -- 0x00000738
    x"00000000", -- 0x0000073c
    x"8fc2000c", -- 0x00000740
    x"00000000", -- 0x00000744
    x"40826000", -- 0x00000748
    x"1000000a", -- 0x0000074c
    x"00000000", -- 0x00000750
    x"8fc2000c", -- 0x00000754
    x"00000000", -- 0x00000758
    x"40826800", -- 0x0000075c
    x"10000005", -- 0x00000760
    x"00000000", -- 0x00000764
    x"8fc2000c", -- 0x00000768
    x"00000000", -- 0x0000076c
    x"40827000", -- 0x00000770
    x"00000000", -- 0x00000774
    x"00000000", -- 0x00000778
    x"03c0e825", -- 0x0000077c
    x"8fbe0004", -- 0x00000780
    x"27bd0008", -- 0x00000784
    x"03e00008", -- 0x00000788
    x"00000000", -- 0x0000078c
    x"27bdffe0", -- 0x00000790
    x"afbf001c", -- 0x00000794
    x"afbe0018", -- 0x00000798
    x"03a0f025", -- 0x0000079c
    x"afc40020", -- 0x000007a0
    x"afc00010", -- 0x000007a4
    x"8fc20020", -- 0x000007a8
    x"00000000", -- 0x000007ac
    x"8c42001c", -- 0x000007b0
    x"00000000", -- 0x000007b4
    x"00021900", -- 0x000007b8
    x"8fc20020", -- 0x000007bc
    x"00000000", -- 0x000007c0
    x"8c420018", -- 0x000007c4
    x"00000000", -- 0x000007c8
    x"000210c0", -- 0x000007cc
    x"00621825", -- 0x000007d0
    x"8fc20020", -- 0x000007d4
    x"00000000", -- 0x000007d8
    x"8c420014", -- 0x000007dc
    x"00000000", -- 0x000007e0
    x"00021080", -- 0x000007e4
    x"00621825", -- 0x000007e8
    x"8fc20020", -- 0x000007ec
    x"00000000", -- 0x000007f0
    x"8c420010", -- 0x000007f4
    x"00000000", -- 0x000007f8
    x"00621025", -- 0x000007fc
    x"8fc30010", -- 0x00000800
    x"00000000", -- 0x00000804
    x"00621025", -- 0x00000808
    x"afc20010", -- 0x0000080c
    x"8fc20020", -- 0x00000810
    x"00000000", -- 0x00000814
    x"8c430000", -- 0x00000818
    x"24020001", -- 0x0000081c
    x"14620022", -- 0x00000820
    x"00000000", -- 0x00000824
    x"8fc20020", -- 0x00000828
    x"00000000", -- 0x0000082c
    x"8c420004", -- 0x00000830
    x"00000000", -- 0x00000834
    x"00402825", -- 0x00000838
    x"3c040003", -- 0x0000083c
    x"0c00012b", -- 0x00000840
    x"00000000", -- 0x00000844
    x"8fc20020", -- 0x00000848
    x"00000000", -- 0x0000084c
    x"8c420008", -- 0x00000850
    x"00000000", -- 0x00000854
    x"00402825", -- 0x00000858
    x"3c020003", -- 0x0000085c
    x"34440004", -- 0x00000860
    x"0c00012b", -- 0x00000864
    x"00000000", -- 0x00000868
    x"8fc20020", -- 0x0000086c
    x"00000000", -- 0x00000870
    x"8c42000c", -- 0x00000874
    x"00000000", -- 0x00000878
    x"00402825", -- 0x0000087c
    x"3c020003", -- 0x00000880
    x"34440008", -- 0x00000884
    x"0c00012b", -- 0x00000888
    x"00000000", -- 0x0000088c
    x"8fc50010", -- 0x00000890
    x"3c020003", -- 0x00000894
    x"3444000c", -- 0x00000898
    x"0c00012b", -- 0x0000089c
    x"00000000", -- 0x000008a0
    x"10000077", -- 0x000008a4
    x"00000000", -- 0x000008a8
    x"8fc20020", -- 0x000008ac
    x"00000000", -- 0x000008b0
    x"8c430000", -- 0x000008b4
    x"24020002", -- 0x000008b8
    x"14620023", -- 0x000008bc
    x"00000000", -- 0x000008c0
    x"8fc20020", -- 0x000008c4
    x"00000000", -- 0x000008c8
    x"8c420004", -- 0x000008cc
    x"00000000", -- 0x000008d0
    x"00402825", -- 0x000008d4
    x"3c020003", -- 0x000008d8
    x"34440010", -- 0x000008dc
    x"0c00012b", -- 0x000008e0
    x"00000000", -- 0x000008e4
    x"8fc20020", -- 0x000008e8
    x"00000000", -- 0x000008ec
    x"8c420008", -- 0x000008f0
    x"00000000", -- 0x000008f4
    x"00402825", -- 0x000008f8
    x"3c020003", -- 0x000008fc
    x"34440014", -- 0x00000900
    x"0c00012b", -- 0x00000904
    x"00000000", -- 0x00000908
    x"8fc20020", -- 0x0000090c
    x"00000000", -- 0x00000910
    x"8c42000c", -- 0x00000914
    x"00000000", -- 0x00000918
    x"00402825", -- 0x0000091c
    x"3c020003", -- 0x00000920
    x"34440018", -- 0x00000924
    x"0c00012b", -- 0x00000928
    x"00000000", -- 0x0000092c
    x"8fc50010", -- 0x00000930
    x"3c020003", -- 0x00000934
    x"3444001c", -- 0x00000938
    x"0c00012b", -- 0x0000093c
    x"00000000", -- 0x00000940
    x"1000004f", -- 0x00000944
    x"00000000", -- 0x00000948
    x"8fc20020", -- 0x0000094c
    x"00000000", -- 0x00000950
    x"8c430000", -- 0x00000954
    x"24020004", -- 0x00000958
    x"14620023", -- 0x0000095c
    x"00000000", -- 0x00000960
    x"8fc20020", -- 0x00000964
    x"00000000", -- 0x00000968
    x"8c420004", -- 0x0000096c
    x"00000000", -- 0x00000970
    x"00402825", -- 0x00000974
    x"3c020003", -- 0x00000978
    x"34440020", -- 0x0000097c
    x"0c00012b", -- 0x00000980
    x"00000000", -- 0x00000984
    x"8fc20020", -- 0x00000988
    x"00000000", -- 0x0000098c
    x"8c420008", -- 0x00000990
    x"00000000", -- 0x00000994
    x"00402825", -- 0x00000998
    x"3c020003", -- 0x0000099c
    x"34440024", -- 0x000009a0
    x"0c00012b", -- 0x000009a4
    x"00000000", -- 0x000009a8
    x"8fc20020", -- 0x000009ac
    x"00000000", -- 0x000009b0
    x"8c42000c", -- 0x000009b4
    x"00000000", -- 0x000009b8
    x"00402825", -- 0x000009bc
    x"3c020003", -- 0x000009c0
    x"34440028", -- 0x000009c4
    x"0c00012b", -- 0x000009c8
    x"00000000", -- 0x000009cc
    x"8fc50010", -- 0x000009d0
    x"3c020003", -- 0x000009d4
    x"3444002c", -- 0x000009d8
    x"0c00012b", -- 0x000009dc
    x"00000000", -- 0x000009e0
    x"10000027", -- 0x000009e4
    x"00000000", -- 0x000009e8
    x"8fc20020", -- 0x000009ec
    x"00000000", -- 0x000009f0
    x"8c430000", -- 0x000009f4
    x"24020008", -- 0x000009f8
    x"14620021", -- 0x000009fc
    x"00000000", -- 0x00000a00
    x"8fc20020", -- 0x00000a04
    x"00000000", -- 0x00000a08
    x"8c420004", -- 0x00000a0c
    x"00000000", -- 0x00000a10
    x"00402825", -- 0x00000a14
    x"3c020003", -- 0x00000a18
    x"34440030", -- 0x00000a1c
    x"0c00012b", -- 0x00000a20
    x"00000000", -- 0x00000a24
    x"8fc20020", -- 0x00000a28
    x"00000000", -- 0x00000a2c
    x"8c420008", -- 0x00000a30
    x"00000000", -- 0x00000a34
    x"00402825", -- 0x00000a38
    x"3c020003", -- 0x00000a3c
    x"34440034", -- 0x00000a40
    x"0c00012b", -- 0x00000a44
    x"00000000", -- 0x00000a48
    x"8fc20020", -- 0x00000a4c
    x"00000000", -- 0x00000a50
    x"8c42000c", -- 0x00000a54
    x"00000000", -- 0x00000a58
    x"00402825", -- 0x00000a5c
    x"3c020003", -- 0x00000a60
    x"34440038", -- 0x00000a64
    x"0c00012b", -- 0x00000a68
    x"00000000", -- 0x00000a6c
    x"8fc50010", -- 0x00000a70
    x"3c020003", -- 0x00000a74
    x"3444003c", -- 0x00000a78
    x"0c00012b", -- 0x00000a7c
    x"00000000", -- 0x00000a80
    x"24040400", -- 0x00000a84
    x"0c00016a", -- 0x00000a88
    x"00000000", -- 0x00000a8c
    x"00000000", -- 0x00000a90
    x"03c0e825", -- 0x00000a94
    x"8fbf001c", -- 0x00000a98
    x"8fbe0018", -- 0x00000a9c
    x"27bd0020", -- 0x00000aa0
    x"03e00008", -- 0x00000aa4
    x"00000000", -- 0x00000aa8
    x"27bdffe8", -- 0x00000aac
    x"afbf0014", -- 0x00000ab0
    x"afbe0010", -- 0x00000ab4
    x"03a0f025", -- 0x00000ab8
    x"afc40018", -- 0x00000abc
    x"8fc20018", -- 0x00000ac0
    x"00000000", -- 0x00000ac4
    x"8c430000", -- 0x00000ac8
    x"24020001", -- 0x00000acc
    x"1462000d", -- 0x00000ad0
    x"00000000", -- 0x00000ad4
    x"8fc20018", -- 0x00000ad8
    x"00000000", -- 0x00000adc
    x"8c420020", -- 0x00000ae0
    x"00000000", -- 0x00000ae4
    x"34420100", -- 0x00000ae8
    x"00402825", -- 0x00000aec
    x"3c020003", -- 0x00000af0
    x"3444000c", -- 0x00000af4
    x"0c00012b", -- 0x00000af8
    x"00000000", -- 0x00000afc
    x"10000035", -- 0x00000b00
    x"00000000", -- 0x00000b04
    x"8fc20018", -- 0x00000b08
    x"00000000", -- 0x00000b0c
    x"8c430000", -- 0x00000b10
    x"24020002", -- 0x00000b14
    x"1462000d", -- 0x00000b18
    x"00000000", -- 0x00000b1c
    x"8fc20018", -- 0x00000b20
    x"00000000", -- 0x00000b24
    x"8c420020", -- 0x00000b28
    x"00000000", -- 0x00000b2c
    x"34420100", -- 0x00000b30
    x"00402825", -- 0x00000b34
    x"3c020003", -- 0x00000b38
    x"3444001c", -- 0x00000b3c
    x"0c00012b", -- 0x00000b40
    x"00000000", -- 0x00000b44
    x"10000023", -- 0x00000b48
    x"00000000", -- 0x00000b4c
    x"8fc20018", -- 0x00000b50
    x"00000000", -- 0x00000b54
    x"8c430000", -- 0x00000b58
    x"24020004", -- 0x00000b5c
    x"1462000d", -- 0x00000b60
    x"00000000", -- 0x00000b64
    x"8fc20018", -- 0x00000b68
    x"00000000", -- 0x00000b6c
    x"8c420020", -- 0x00000b70
    x"00000000", -- 0x00000b74
    x"34420100", -- 0x00000b78
    x"00402825", -- 0x00000b7c
    x"3c020003", -- 0x00000b80
    x"3444002c", -- 0x00000b84
    x"0c00012b", -- 0x00000b88
    x"00000000", -- 0x00000b8c
    x"10000011", -- 0x00000b90
    x"00000000", -- 0x00000b94
    x"8fc20018", -- 0x00000b98
    x"00000000", -- 0x00000b9c
    x"8c430000", -- 0x00000ba0
    x"24020008", -- 0x00000ba4
    x"1462000b", -- 0x00000ba8
    x"00000000", -- 0x00000bac
    x"8fc20018", -- 0x00000bb0
    x"00000000", -- 0x00000bb4
    x"8c420020", -- 0x00000bb8
    x"00000000", -- 0x00000bbc
    x"34420100", -- 0x00000bc0
    x"00402825", -- 0x00000bc4
    x"3c020003", -- 0x00000bc8
    x"3444003c", -- 0x00000bcc
    x"0c00012b", -- 0x00000bd0
    x"00000000", -- 0x00000bd4
    x"00000000", -- 0x00000bd8
    x"03c0e825", -- 0x00000bdc
    x"8fbf0014", -- 0x00000be0
    x"8fbe0010", -- 0x00000be4
    x"27bd0018", -- 0x00000be8
    x"03e00008", -- 0x00000bec
    x"00000000", -- 0x00000bf0
    x"27bdffe8", -- 0x00000bf4
    x"afbf0014", -- 0x00000bf8
    x"afbe0010", -- 0x00000bfc
    x"03a0f025", -- 0x00000c00
    x"afc40018", -- 0x00000c04
    x"8fc20018", -- 0x00000c08
    x"00000000", -- 0x00000c0c
    x"8c430000", -- 0x00000c10
    x"24020001", -- 0x00000c14
    x"1462000d", -- 0x00000c18
    x"00000000", -- 0x00000c1c
    x"8fc20018", -- 0x00000c20
    x"00000000", -- 0x00000c24
    x"8c420020", -- 0x00000c28
    x"00000000", -- 0x00000c2c
    x"34420200", -- 0x00000c30
    x"00402825", -- 0x00000c34
    x"3c020003", -- 0x00000c38
    x"3444000c", -- 0x00000c3c
    x"0c00012b", -- 0x00000c40
    x"00000000", -- 0x00000c44
    x"10000035", -- 0x00000c48
    x"00000000", -- 0x00000c4c
    x"8fc20018", -- 0x00000c50
    x"00000000", -- 0x00000c54
    x"8c430000", -- 0x00000c58
    x"24020002", -- 0x00000c5c
    x"1462000d", -- 0x00000c60
    x"00000000", -- 0x00000c64
    x"8fc20018", -- 0x00000c68
    x"00000000", -- 0x00000c6c
    x"8c420020", -- 0x00000c70
    x"00000000", -- 0x00000c74
    x"34420200", -- 0x00000c78
    x"00402825", -- 0x00000c7c
    x"3c020003", -- 0x00000c80
    x"3444001c", -- 0x00000c84
    x"0c00012b", -- 0x00000c88
    x"00000000", -- 0x00000c8c
    x"10000023", -- 0x00000c90
    x"00000000", -- 0x00000c94
    x"8fc20018", -- 0x00000c98
    x"00000000", -- 0x00000c9c
    x"8c430000", -- 0x00000ca0
    x"24020004", -- 0x00000ca4
    x"1462000d", -- 0x00000ca8
    x"00000000", -- 0x00000cac
    x"8fc20018", -- 0x00000cb0
    x"00000000", -- 0x00000cb4
    x"8c420020", -- 0x00000cb8
    x"00000000", -- 0x00000cbc
    x"34420200", -- 0x00000cc0
    x"00402825", -- 0x00000cc4
    x"3c020003", -- 0x00000cc8
    x"3444002c", -- 0x00000ccc
    x"0c00012b", -- 0x00000cd0
    x"00000000", -- 0x00000cd4
    x"10000011", -- 0x00000cd8
    x"00000000", -- 0x00000cdc
    x"8fc20018", -- 0x00000ce0
    x"00000000", -- 0x00000ce4
    x"8c430000", -- 0x00000ce8
    x"24020008", -- 0x00000cec
    x"1462000b", -- 0x00000cf0
    x"00000000", -- 0x00000cf4
    x"8fc20018", -- 0x00000cf8
    x"00000000", -- 0x00000cfc
    x"8c420020", -- 0x00000d00
    x"00000000", -- 0x00000d04
    x"34420200", -- 0x00000d08
    x"00402825", -- 0x00000d0c
    x"3c020003", -- 0x00000d10
    x"3444003c", -- 0x00000d14
    x"0c00012b", -- 0x00000d18
    x"00000000", -- 0x00000d1c
    x"00000000", -- 0x00000d20
    x"03c0e825", -- 0x00000d24
    x"8fbf0014", -- 0x00000d28
    x"8fbe0010", -- 0x00000d2c
    x"27bd0018", -- 0x00000d30
    x"03e00008", -- 0x00000d34
    x"00000000", -- 0x00000d38
    x"27bdfff8", -- 0x00000d3c
    x"afbe0004", -- 0x00000d40
    x"03a0f025", -- 0x00000d44
    x"afc40008", -- 0x00000d48
    x"00000000", -- 0x00000d4c
    x"03c0e825", -- 0x00000d50
    x"8fbe0004", -- 0x00000d54
    x"27bd0008", -- 0x00000d58
    x"03e00008", -- 0x00000d5c
    x"00000000", -- 0x00000d60
    x"27bdfff8", -- 0x00000d64
    x"afbe0004", -- 0x00000d68
    x"03a0f025", -- 0x00000d6c
    x"2402ffff", -- 0x00000d70
    x"03c0e825", -- 0x00000d74
    x"8fbe0004", -- 0x00000d78
    x"27bd0008", -- 0x00000d7c
    x"03e00008", -- 0x00000d80
    x"00000000", -- 0x00000d84
    x"27bdffe0", -- 0x00000d88
    x"afbf001c", -- 0x00000d8c
    x"afbe0018", -- 0x00000d90
    x"03a0f025", -- 0x00000d94
    x"3c020003", -- 0x00000d98
    x"34440040", -- 0x00000d9c
    x"0c00013a", -- 0x00000da0
    x"00000000", -- 0x00000da4
    x"afc20010", -- 0x00000da8
    x"8fc30010", -- 0x00000dac
    x"3c020001", -- 0x00000db0
    x"00621024", -- 0x00000db4
    x"10400026", -- 0x00000db8
    x"00000000", -- 0x00000dbc
    x"8f83008c", -- 0x00000dc0
    x"8f820000", -- 0x00000dc4
    x"00000000", -- 0x00000dc8
    x"00621021", -- 0x00000dcc
    x"00402825", -- 0x00000dd0
    x"3c020003", -- 0x00000dd4
    x"34440014", -- 0x00000dd8
    x"0c00012b", -- 0x00000ddc
    x"00000000", -- 0x00000de0
    x"8f820084", -- 0x00000de4
    x"00000000", -- 0x00000de8
    x"00402025", -- 0x00000dec
    x"0c0002ab", -- 0x00000df0
    x"00000000", -- 0x00000df4
    x"8f820088", -- 0x00000df8
    x"00000000", -- 0x00000dfc
    x"00402025", -- 0x00000e00
    x"0c0002fd", -- 0x00000e04
    x"00000000", -- 0x00000e08
    x"8f820088", -- 0x00000e0c
    x"00000000", -- 0x00000e10
    x"00402025", -- 0x00000e14
    x"0c0002ab", -- 0x00000e18
    x"00000000", -- 0x00000e1c
    x"8f820000", -- 0x00000e20
    x"00000000", -- 0x00000e24
    x"24420040", -- 0x00000e28
    x"2c420400", -- 0x00000e2c
    x"14400004", -- 0x00000e30
    x"00000000", -- 0x00000e34
    x"af800000", -- 0x00000e38
    x"10000005", -- 0x00000e3c
    x"00000000", -- 0x00000e40
    x"8f820000", -- 0x00000e44
    x"00000000", -- 0x00000e48
    x"24420040", -- 0x00000e4c
    x"af820000", -- 0x00000e50
    x"8fc30010", -- 0x00000e54
    x"3c020002", -- 0x00000e58
    x"00621024", -- 0x00000e5c
    x"10400021", -- 0x00000e60
    x"00000000", -- 0x00000e64
    x"8f820084", -- 0x00000e68
    x"00000000", -- 0x00000e6c
    x"00402025", -- 0x00000e70
    x"0c0002fd", -- 0x00000e74
    x"00000000", -- 0x00000e78
    x"8f83008c", -- 0x00000e7c
    x"8f820004", -- 0x00000e80
    x"00000000", -- 0x00000e84
    x"00621021", -- 0x00000e88
    x"00402825", -- 0x00000e8c
    x"3c020003", -- 0x00000e90
    x"34440020", -- 0x00000e94
    x"0c00012b", -- 0x00000e98
    x"00000000", -- 0x00000e9c
    x"8f820080", -- 0x00000ea0
    x"00000000", -- 0x00000ea4
    x"00402025", -- 0x00000ea8
    x"0c0002ab", -- 0x00000eac
    x"00000000", -- 0x00000eb0
    x"8f820004", -- 0x00000eb4
    x"00000000", -- 0x00000eb8
    x"24420040", -- 0x00000ebc
    x"2c420400", -- 0x00000ec0
    x"14400004", -- 0x00000ec4
    x"00000000", -- 0x00000ec8
    x"af800004", -- 0x00000ecc
    x"10000005", -- 0x00000ed0
    x"00000000", -- 0x00000ed4
    x"8f820004", -- 0x00000ed8
    x"00000000", -- 0x00000edc
    x"24420040", -- 0x00000ee0
    x"af820004", -- 0x00000ee4
    x"8fc30010", -- 0x00000ee8
    x"3c020004", -- 0x00000eec
    x"00621024", -- 0x00000ef0
    x"10400006", -- 0x00000ef4
    x"00000000", -- 0x00000ef8
    x"8f820080", -- 0x00000efc
    x"00000000", -- 0x00000f00
    x"00402025", -- 0x00000f04
    x"0c0002fd", -- 0x00000f08
    x"00000000", -- 0x00000f0c
    x"00000000", -- 0x00000f10
    x"03c0e825", -- 0x00000f14
    x"8fbf001c", -- 0x00000f18
    x"8fbe0018", -- 0x00000f1c
    x"27bd0020", -- 0x00000f20
    x"03e00008", -- 0x00000f24
    x"00000000", -- 0x00000f28
    x"27bdfb30", -- 0x00000f2c
    x"afbf04cc", -- 0x00000f30
    x"afbe04c8", -- 0x00000f34
    x"03a0f025", -- 0x00000f38
    x"afa00010", -- 0x00000f3c
    x"00003825", -- 0x00000f40
    x"24060008", -- 0x00000f44
    x"3c020001", -- 0x00000f48
    x"3445c200", -- 0x00000f4c
    x"34048200", -- 0x00000f50
    x"0c00080e", -- 0x00000f54
    x"00000000", -- 0x00000f58
    x"afc0045c", -- 0x00000f5c
    x"afc00460", -- 0x00000f60
    x"afc00464", -- 0x00000f64
    x"afc00468", -- 0x00000f68
    x"afc0046c", -- 0x00000f6c
    x"afc00470", -- 0x00000f70
    x"afc00474", -- 0x00000f74
    x"afc00478", -- 0x00000f78
    x"afc0047c", -- 0x00000f7c
    x"24020001", -- 0x00000f80
    x"afc2045c", -- 0x00000f84
    x"34028204", -- 0x00000f88
    x"afc20460", -- 0x00000f8c
    x"27c2001c", -- 0x00000f90
    x"afc20464", -- 0x00000f94
    x"24020040", -- 0x00000f98
    x"afc20468", -- 0x00000f9c
    x"24020001", -- 0x00000fa0
    x"afc2046c", -- 0x00000fa4
    x"24020001", -- 0x00000fa8
    x"afc20470", -- 0x00000fac
    x"24020001", -- 0x00000fb0
    x"afc20474", -- 0x00000fb4
    x"24020001", -- 0x00000fb8
    x"afc20478", -- 0x00000fbc
    x"27c2045c", -- 0x00000fc0
    x"af820088", -- 0x00000fc4
    x"afc00480", -- 0x00000fc8
    x"afc00484", -- 0x00000fcc
    x"afc00488", -- 0x00000fd0
    x"afc0048c", -- 0x00000fd4
    x"afc00490", -- 0x00000fd8
    x"afc00494", -- 0x00000fdc
    x"afc00498", -- 0x00000fe0
    x"afc0049c", -- 0x00000fe4
    x"afc004a0", -- 0x00000fe8
    x"24020002", -- 0x00000fec
    x"afc20480", -- 0x00000ff0
    x"27c2001c", -- 0x00000ff4
    x"afc20484", -- 0x00000ff8
    x"24020040", -- 0x00000ffc
    x"afc2048c", -- 0x00001000
    x"24020001", -- 0x00001004
    x"afc20498", -- 0x00001008
    x"27c20480", -- 0x0000100c
    x"af820084", -- 0x00001010
    x"afc004a4", -- 0x00001014
    x"afc004a8", -- 0x00001018
    x"afc004ac", -- 0x0000101c
    x"afc004b0", -- 0x00001020
    x"afc004b4", -- 0x00001024
    x"afc004b8", -- 0x00001028
    x"afc004bc", -- 0x0000102c
    x"afc004c0", -- 0x00001030
    x"afc004c4", -- 0x00001034
    x"24020004", -- 0x00001038
    x"afc204a4", -- 0x0000103c
    x"34028200", -- 0x00001040
    x"afc204ac", -- 0x00001044
    x"24020040", -- 0x00001048
    x"afc204b0", -- 0x0000104c
    x"24020002", -- 0x00001050
    x"afc204b4", -- 0x00001054
    x"24020001", -- 0x00001058
    x"afc204b8", -- 0x0000105c
    x"24020001", -- 0x00001060
    x"afc204bc", -- 0x00001064
    x"24020001", -- 0x00001068
    x"afc204c0", -- 0x0000106c
    x"27c204a4", -- 0x00001070
    x"af820080", -- 0x00001074
    x"27c2045c", -- 0x00001078
    x"00402025", -- 0x0000107c
    x"0c0001e4", -- 0x00001080
    x"00000000", -- 0x00001084
    x"27c20480", -- 0x00001088
    x"00402025", -- 0x0000108c
    x"0c0001e4", -- 0x00001090
    x"00000000", -- 0x00001094
    x"27c204a4", -- 0x00001098
    x"00402025", -- 0x0000109c
    x"0c0001e4", -- 0x000010a0
    x"00000000", -- 0x000010a4
    x"27c2005c", -- 0x000010a8
    x"af82008c", -- 0x000010ac
    x"34048208", -- 0x000010b0
    x"0c00013a", -- 0x000010b4
    x"00000000", -- 0x000010b8
    x"00401825", -- 0x000010bc
    x"3c020200", -- 0x000010c0
    x"00621025", -- 0x000010c4
    x"00402825", -- 0x000010c8
    x"34048208", -- 0x000010cc
    x"0c00012b", -- 0x000010d0
    x"00000000", -- 0x000010d4
    x"3c020003", -- 0x000010d8
    x"3444000c", -- 0x000010dc
    x"0c00013a", -- 0x000010e0
    x"00000000", -- 0x000010e4
    x"afc2047c", -- 0x000010e8
    x"3c020003", -- 0x000010ec
    x"3444001c", -- 0x000010f0
    x"0c00013a", -- 0x000010f4
    x"00000000", -- 0x000010f8
    x"afc204a0", -- 0x000010fc
    x"3c020003", -- 0x00001100
    x"3444002c", -- 0x00001104
    x"0c00013a", -- 0x00001108
    x"00000000", -- 0x0000110c
    x"afc204c4", -- 0x00001110
    x"27c2045c", -- 0x00001114
    x"00402025", -- 0x00001118
    x"0c0002ab", -- 0x0000111c
    x"00000000", -- 0x00001120
    x"8fc20018", -- 0x00001124
    x"00000000", -- 0x00001128
    x"24420001", -- 0x0000112c
    x"afc20018", -- 0x00001130
    x"1000fffb", -- 0x00001134
    x"00000000", -- 0x00001138
    x"27bdfff0", -- 0x0000113c
    x"afbe000c", -- 0x00001140
    x"03a0f025", -- 0x00001144
    x"afc40010", -- 0x00001148
    x"afc50014", -- 0x0000114c
    x"afc60018", -- 0x00001150
    x"8fc20010", -- 0x00001154
    x"00000000", -- 0x00001158
    x"afc20000", -- 0x0000115c
    x"8fc20014", -- 0x00001160
    x"00000000", -- 0x00001164
    x"afc20004", -- 0x00001168
    x"1000000c", -- 0x0000116c
    x"00000000", -- 0x00001170
    x"8fc20000", -- 0x00001174
    x"00000000", -- 0x00001178
    x"24430001", -- 0x0000117c
    x"afc30000", -- 0x00001180
    x"8fc30004", -- 0x00001184
    x"00000000", -- 0x00001188
    x"24640001", -- 0x0000118c
    x"afc40004", -- 0x00001190
    x"90630000", -- 0x00001194
    x"00000000", -- 0x00001198
    x"a0430000", -- 0x0000119c
    x"8fc20018", -- 0x000011a0
    x"00000000", -- 0x000011a4
    x"2443ffff", -- 0x000011a8
    x"afc30018", -- 0x000011ac
    x"1440fff0", -- 0x000011b0
    x"00000000", -- 0x000011b4
    x"8fc20010", -- 0x000011b8
    x"03c0e825", -- 0x000011bc
    x"8fbe000c", -- 0x000011c0
    x"27bd0010", -- 0x000011c4
    x"03e00008", -- 0x000011c8
    x"00000000", -- 0x000011cc
    x"27bdfff0", -- 0x000011d0
    x"afbe000c", -- 0x000011d4
    x"03a0f025", -- 0x000011d8
    x"afc40010", -- 0x000011dc
    x"afc50014", -- 0x000011e0
    x"afc60018", -- 0x000011e4
    x"8fc20010", -- 0x000011e8
    x"00000000", -- 0x000011ec
    x"afc20000", -- 0x000011f0
    x"10000009", -- 0x000011f4
    x"00000000", -- 0x000011f8
    x"8fc20000", -- 0x000011fc
    x"00000000", -- 0x00001200
    x"24430001", -- 0x00001204
    x"afc30000", -- 0x00001208
    x"8fc30014", -- 0x0000120c
    x"00000000", -- 0x00001210
    x"306300ff", -- 0x00001214
    x"a0430000", -- 0x00001218
    x"8fc20018", -- 0x0000121c
    x"00000000", -- 0x00001220
    x"2443ffff", -- 0x00001224
    x"afc30018", -- 0x00001228
    x"1440fff3", -- 0x0000122c
    x"00000000", -- 0x00001230
    x"8fc20010", -- 0x00001234
    x"03c0e825", -- 0x00001238
    x"8fbe000c", -- 0x0000123c
    x"27bd0010", -- 0x00001240
    x"03e00008", -- 0x00001244
    x"00000000", -- 0x00001248
    x"27bdffe8", -- 0x0000124c
    x"afbf0014", -- 0x00001250
    x"afbe0010", -- 0x00001254
    x"03a0f025", -- 0x00001258
    x"27830000", -- 0x0000125c
    x"2782e207", -- 0x00001260
    x"10620009", -- 0x00001264
    x"00000000", -- 0x00001268
    x"27830000", -- 0x0000126c
    x"27820000", -- 0x00001270
    x"00621023", -- 0x00001274
    x"00403025", -- 0x00001278
    x"2785e207", -- 0x0000127c
    x"27840000", -- 0x00001280
    x"0c00044f", -- 0x00001284
    x"00000000", -- 0x00001288
    x"27830080", -- 0x0000128c
    x"27820000", -- 0x00001290
    x"00621023", -- 0x00001294
    x"00403025", -- 0x00001298
    x"00002825", -- 0x0000129c
    x"27840000", -- 0x000012a0
    x"0c000474", -- 0x000012a4
    x"00000000", -- 0x000012a8
    x"0c0003cb", -- 0x000012ac
    x"00000000", -- 0x000012b0
    x"1000ffff", -- 0x000012b4
    x"00000000", -- 0x000012b8
    x"27bdffe8", -- 0x000012bc
    x"afbf0014", -- 0x000012c0
    x"afbe0010", -- 0x000012c4
    x"03a0f025", -- 0x000012c8
    x"afc40018", -- 0x000012cc
    x"1000000a", -- 0x000012d0
    x"00000000", -- 0x000012d4
    x"8fc20018", -- 0x000012d8
    x"00000000", -- 0x000012dc
    x"24430001", -- 0x000012e0
    x"afc30018", -- 0x000012e4
    x"90420000", -- 0x000012e8
    x"00000000", -- 0x000012ec
    x"00402025", -- 0x000012f0
    x"0c000856", -- 0x000012f4
    x"00000000", -- 0x000012f8
    x"8fc20018", -- 0x000012fc
    x"00000000", -- 0x00001300
    x"90420000", -- 0x00001304
    x"00000000", -- 0x00001308
    x"1440fff2", -- 0x0000130c
    x"00000000", -- 0x00001310
    x"2404000a", -- 0x00001314
    x"0c000856", -- 0x00001318
    x"00000000", -- 0x0000131c
    x"00001025", -- 0x00001320
    x"03c0e825", -- 0x00001324
    x"8fbf0014", -- 0x00001328
    x"8fbe0010", -- 0x0000132c
    x"27bd0018", -- 0x00001330
    x"03e00008", -- 0x00001334
    x"00000000", -- 0x00001338
    x"27bdffe8", -- 0x0000133c
    x"afbf0014", -- 0x00001340
    x"afbe0010", -- 0x00001344
    x"03a0f025", -- 0x00001348
    x"afc40018", -- 0x0000134c
    x"afc5001c", -- 0x00001350
    x"8fc20018", -- 0x00001354
    x"00000000", -- 0x00001358
    x"10400012", -- 0x0000135c
    x"00000000", -- 0x00001360
    x"8fc20018", -- 0x00001364
    x"00000000", -- 0x00001368
    x"8c420000", -- 0x0000136c
    x"8fc3001c", -- 0x00001370
    x"00000000", -- 0x00001374
    x"306300ff", -- 0x00001378
    x"a0430000", -- 0x0000137c
    x"8fc20018", -- 0x00001380
    x"00000000", -- 0x00001384
    x"8c420000", -- 0x00001388
    x"00000000", -- 0x0000138c
    x"24430001", -- 0x00001390
    x"8fc20018", -- 0x00001394
    x"00000000", -- 0x00001398
    x"ac430000", -- 0x0000139c
    x"10000004", -- 0x000013a0
    x"00000000", -- 0x000013a4
    x"8fc4001c", -- 0x000013a8
    x"0c000856", -- 0x000013ac
    x"00000000", -- 0x000013b0
    x"00000000", -- 0x000013b4
    x"03c0e825", -- 0x000013b8
    x"8fbf0014", -- 0x000013bc
    x"8fbe0010", -- 0x000013c0
    x"27bd0018", -- 0x000013c4
    x"03e00008", -- 0x000013c8
    x"00000000", -- 0x000013cc
    x"27bdffd8", -- 0x000013d0
    x"afbf0024", -- 0x000013d4
    x"afbe0020", -- 0x000013d8
    x"afb3001c", -- 0x000013dc
    x"afb20018", -- 0x000013e0
    x"afb10014", -- 0x000013e4
    x"afb00010", -- 0x000013e8
    x"03a0f025", -- 0x000013ec
    x"afc40028", -- 0x000013f0
    x"afc5002c", -- 0x000013f4
    x"afc60030", -- 0x000013f8
    x"afc70034", -- 0x000013fc
    x"00008025", -- 0x00001400
    x"24130020", -- 0x00001404
    x"8fc20030", -- 0x00001408
    x"00000000", -- 0x0000140c
    x"1840001d", -- 0x00001410
    x"00000000", -- 0x00001414
    x"00008825", -- 0x00001418
    x"8fd2002c", -- 0x0000141c
    x"10000003", -- 0x00001420
    x"00000000", -- 0x00001424
    x"26310001", -- 0x00001428
    x"26520001", -- 0x0000142c
    x"92420000", -- 0x00001430
    x"00000000", -- 0x00001434
    x"1440fffb", -- 0x00001438
    x"00000000", -- 0x0000143c
    x"8fc20030", -- 0x00001440
    x"00000000", -- 0x00001444
    x"0222102a", -- 0x00001448
    x"14400004", -- 0x0000144c
    x"00000000", -- 0x00001450
    x"afc00030", -- 0x00001454
    x"10000005", -- 0x00001458
    x"00000000", -- 0x0000145c
    x"8fc20030", -- 0x00001460
    x"00000000", -- 0x00001464
    x"00511023", -- 0x00001468
    x"afc20030", -- 0x0000146c
    x"8fc20034", -- 0x00001470
    x"00000000", -- 0x00001474
    x"30420002", -- 0x00001478
    x"10400002", -- 0x0000147c
    x"00000000", -- 0x00001480
    x"24130030", -- 0x00001484
    x"8fc20034", -- 0x00001488
    x"00000000", -- 0x0000148c
    x"30420001", -- 0x00001490
    x"1440001f", -- 0x00001494
    x"00000000", -- 0x00001498
    x"1000000a", -- 0x0000149c
    x"00000000", -- 0x000014a0
    x"02602825", -- 0x000014a4
    x"8fc40028", -- 0x000014a8
    x"0c0004cf", -- 0x000014ac
    x"00000000", -- 0x000014b0
    x"26100001", -- 0x000014b4
    x"8fc20030", -- 0x000014b8
    x"00000000", -- 0x000014bc
    x"2442ffff", -- 0x000014c0
    x"afc20030", -- 0x000014c4
    x"8fc20030", -- 0x000014c8
    x"00000000", -- 0x000014cc
    x"1c40fff4", -- 0x000014d0
    x"00000000", -- 0x000014d4
    x"1000000e", -- 0x000014d8
    x"00000000", -- 0x000014dc
    x"8fc2002c", -- 0x000014e0
    x"00000000", -- 0x000014e4
    x"90420000", -- 0x000014e8
    x"00000000", -- 0x000014ec
    x"00402825", -- 0x000014f0
    x"8fc40028", -- 0x000014f4
    x"0c0004cf", -- 0x000014f8
    x"00000000", -- 0x000014fc
    x"26100001", -- 0x00001500
    x"8fc2002c", -- 0x00001504
    x"00000000", -- 0x00001508
    x"24420001", -- 0x0000150c
    x"afc2002c", -- 0x00001510
    x"8fc2002c", -- 0x00001514
    x"00000000", -- 0x00001518
    x"90420000", -- 0x0000151c
    x"00000000", -- 0x00001520
    x"1440ffee", -- 0x00001524
    x"00000000", -- 0x00001528
    x"1000000a", -- 0x0000152c
    x"00000000", -- 0x00001530
    x"02602825", -- 0x00001534
    x"8fc40028", -- 0x00001538
    x"0c0004cf", -- 0x0000153c
    x"00000000", -- 0x00001540
    x"26100001", -- 0x00001544
    x"8fc20030", -- 0x00001548
    x"00000000", -- 0x0000154c
    x"2442ffff", -- 0x00001550
    x"afc20030", -- 0x00001554
    x"8fc20030", -- 0x00001558
    x"00000000", -- 0x0000155c
    x"1c40fff4", -- 0x00001560
    x"00000000", -- 0x00001564
    x"02001025", -- 0x00001568
    x"03c0e825", -- 0x0000156c
    x"8fbf0024", -- 0x00001570
    x"8fbe0020", -- 0x00001574
    x"8fb3001c", -- 0x00001578
    x"8fb20018", -- 0x0000157c
    x"8fb10014", -- 0x00001580
    x"8fb00010", -- 0x00001584
    x"27bd0028", -- 0x00001588
    x"03e00008", -- 0x0000158c
    x"00000000", -- 0x00001590
    x"27bdffc8", -- 0x00001594
    x"afbf0034", -- 0x00001598
    x"afbe0030", -- 0x0000159c
    x"afb3002c", -- 0x000015a0
    x"afb20028", -- 0x000015a4
    x"afb10024", -- 0x000015a8
    x"afb00020", -- 0x000015ac
    x"03a0f025", -- 0x000015b0
    x"afc40038", -- 0x000015b4
    x"afc5003c", -- 0x000015b8
    x"afc60040", -- 0x000015bc
    x"afc70044", -- 0x000015c0
    x"00009825", -- 0x000015c4
    x"00009025", -- 0x000015c8
    x"8fdf003c", -- 0x000015cc
    x"8fc2003c", -- 0x000015d0
    x"00000000", -- 0x000015d4
    x"1440000d", -- 0x000015d8
    x"00000000", -- 0x000015dc
    x"24020030", -- 0x000015e0
    x"a3c20010", -- 0x000015e4
    x"a3c00011", -- 0x000015e8
    x"8fc7004c", -- 0x000015ec
    x"8fc60048", -- 0x000015f0
    x"27c20010", -- 0x000015f4
    x"00402825", -- 0x000015f8
    x"8fc40038", -- 0x000015fc
    x"0c0004f4", -- 0x00001600
    x"00000000", -- 0x00001604
    x"1000004e", -- 0x00001608
    x"00000000", -- 0x0000160c
    x"8fc20044", -- 0x00001610
    x"00000000", -- 0x00001614
    x"1040000e", -- 0x00001618
    x"00000000", -- 0x0000161c
    x"8fc30040", -- 0x00001620
    x"2402000a", -- 0x00001624
    x"1462000a", -- 0x00001628
    x"00000000", -- 0x0000162c
    x"8fc2003c", -- 0x00001630
    x"00000000", -- 0x00001634
    x"04410006", -- 0x00001638
    x"00000000", -- 0x0000163c
    x"24130001", -- 0x00001640
    x"8fc2003c", -- 0x00001644
    x"00000000", -- 0x00001648
    x"00021023", -- 0x0000164c
    x"0040f825", -- 0x00001650
    x"27d0001b", -- 0x00001654
    x"a2000000", -- 0x00001658
    x"10000017", -- 0x0000165c
    x"00000000", -- 0x00001660
    x"8fc20040", -- 0x00001664
    x"00000000", -- 0x00001668
    x"03e2001b", -- 0x0000166c
    x"00001010", -- 0x00001670
    x"00408825", -- 0x00001674
    x"2a22000a", -- 0x00001678
    x"14400005", -- 0x0000167c
    x"00000000", -- 0x00001680
    x"8fc20050", -- 0x00001684
    x"00000000", -- 0x00001688
    x"2442ffc6", -- 0x0000168c
    x"02228821", -- 0x00001690
    x"2610ffff", -- 0x00001694
    x"322200ff", -- 0x00001698
    x"24420030", -- 0x0000169c
    x"304200ff", -- 0x000016a0
    x"a2020000", -- 0x000016a4
    x"8fc20040", -- 0x000016a8
    x"00000000", -- 0x000016ac
    x"03e2001b", -- 0x000016b0
    x"00001010", -- 0x000016b4
    x"0000f812", -- 0x000016b8
    x"17e0ffe9", -- 0x000016bc
    x"00000000", -- 0x000016c0
    x"12600018", -- 0x000016c4
    x"00000000", -- 0x000016c8
    x"8fc20048", -- 0x000016cc
    x"00000000", -- 0x000016d0
    x"10400011", -- 0x000016d4
    x"00000000", -- 0x000016d8
    x"8fc2004c", -- 0x000016dc
    x"00000000", -- 0x000016e0
    x"30420002", -- 0x000016e4
    x"1040000c", -- 0x000016e8
    x"00000000", -- 0x000016ec
    x"2405002d", -- 0x000016f0
    x"8fc40038", -- 0x000016f4
    x"0c0004cf", -- 0x000016f8
    x"00000000", -- 0x000016fc
    x"26520001", -- 0x00001700
    x"8fc20048", -- 0x00001704
    x"00000000", -- 0x00001708
    x"2442ffff", -- 0x0000170c
    x"afc20048", -- 0x00001710
    x"10000004", -- 0x00001714
    x"00000000", -- 0x00001718
    x"2610ffff", -- 0x0000171c
    x"2402002d", -- 0x00001720
    x"a2020000", -- 0x00001724
    x"8fc7004c", -- 0x00001728
    x"8fc60048", -- 0x0000172c
    x"02002825", -- 0x00001730
    x"8fc40038", -- 0x00001734
    x"0c0004f4", -- 0x00001738
    x"00000000", -- 0x0000173c
    x"00521021", -- 0x00001740
    x"03c0e825", -- 0x00001744
    x"8fbf0034", -- 0x00001748
    x"8fbe0030", -- 0x0000174c
    x"8fb3002c", -- 0x00001750
    x"8fb20028", -- 0x00001754
    x"8fb10024", -- 0x00001758
    x"8fb00020", -- 0x0000175c
    x"27bd0038", -- 0x00001760
    x"03e00008", -- 0x00001764
    x"00000000", -- 0x00001768
    x"27bdffc0", -- 0x0000176c
    x"afbf003c", -- 0x00001770
    x"afbe0038", -- 0x00001774
    x"afb30034", -- 0x00001778
    x"afb20030", -- 0x0000177c
    x"afb1002c", -- 0x00001780
    x"afb00028", -- 0x00001784
    x"03a0f025", -- 0x00001788
    x"afc40040", -- 0x0000178c
    x"afc50044", -- 0x00001790
    x"00008825", -- 0x00001794
    x"8fc20044", -- 0x00001798
    x"00000000", -- 0x0000179c
    x"24430004", -- 0x000017a0
    x"afc30044", -- 0x000017a4
    x"8c420000", -- 0x000017a8
    x"00000000", -- 0x000017ac
    x"00408025", -- 0x000017b0
    x"100000c5", -- 0x000017b4
    x"00000000", -- 0x000017b8
    x"92030000", -- 0x000017bc
    x"24020025", -- 0x000017c0
    x"146200b9", -- 0x000017c4
    x"00000000", -- 0x000017c8
    x"26100001", -- 0x000017cc
    x"00009825", -- 0x000017d0
    x"02609025", -- 0x000017d4
    x"92020000", -- 0x000017d8
    x"00000000", -- 0x000017dc
    x"104000c0", -- 0x000017e0
    x"00000000", -- 0x000017e4
    x"92030000", -- 0x000017e8
    x"24020025", -- 0x000017ec
    x"106200ad", -- 0x000017f0
    x"00000000", -- 0x000017f4
    x"92030000", -- 0x000017f8
    x"2402002d", -- 0x000017fc
    x"14620007", -- 0x00001800
    x"00000000", -- 0x00001804
    x"26100001", -- 0x00001808
    x"24130001", -- 0x0000180c
    x"10000003", -- 0x00001810
    x"00000000", -- 0x00001814
    x"26100001", -- 0x00001818
    x"36730002", -- 0x0000181c
    x"92030000", -- 0x00001820
    x"24020030", -- 0x00001824
    x"1062fffb", -- 0x00001828
    x"00000000", -- 0x0000182c
    x"1000000a", -- 0x00001830
    x"00000000", -- 0x00001834
    x"02401025", -- 0x00001838
    x"00021040", -- 0x0000183c
    x"00021880", -- 0x00001840
    x"00439021", -- 0x00001844
    x"92020000", -- 0x00001848
    x"00000000", -- 0x0000184c
    x"2442ffd0", -- 0x00001850
    x"02429021", -- 0x00001854
    x"26100001", -- 0x00001858
    x"92020000", -- 0x0000185c
    x"00000000", -- 0x00001860
    x"2c420030", -- 0x00001864
    x"14400006", -- 0x00001868
    x"00000000", -- 0x0000186c
    x"92020000", -- 0x00001870
    x"00000000", -- 0x00001874
    x"2c42003a", -- 0x00001878
    x"1440ffee", -- 0x0000187c
    x"00000000", -- 0x00001880
    x"92030000", -- 0x00001884
    x"24020073", -- 0x00001888
    x"14620017", -- 0x0000188c
    x"00000000", -- 0x00001890
    x"8fc20044", -- 0x00001894
    x"00000000", -- 0x00001898
    x"24430004", -- 0x0000189c
    x"afc30044", -- 0x000018a0
    x"8c5f0000", -- 0x000018a4
    x"00000000", -- 0x000018a8
    x"13e00004", -- 0x000018ac
    x"00000000", -- 0x000018b0
    x"03e01025", -- 0x000018b4
    x"10000003", -- 0x000018b8
    x"00000000", -- 0x000018bc
    x"3c020000", -- 0x000018c0
    x"24422200", -- 0x000018c4
    x"02603825", -- 0x000018c8
    x"02403025", -- 0x000018cc
    x"00402825", -- 0x000018d0
    x"8fc40040", -- 0x000018d4
    x"0c0004f4", -- 0x000018d8
    x"00000000", -- 0x000018dc
    x"02228821", -- 0x000018e0
    x"10000078", -- 0x000018e4
    x"00000000", -- 0x000018e8
    x"92030000", -- 0x000018ec
    x"24020064", -- 0x000018f0
    x"14620013", -- 0x000018f4
    x"00000000", -- 0x000018f8
    x"8fc20044", -- 0x000018fc
    x"00000000", -- 0x00001900
    x"24430004", -- 0x00001904
    x"afc30044", -- 0x00001908
    x"8c430000", -- 0x0000190c
    x"24020061", -- 0x00001910
    x"afa20018", -- 0x00001914
    x"afb30014", -- 0x00001918
    x"afb20010", -- 0x0000191c
    x"24070001", -- 0x00001920
    x"2406000a", -- 0x00001924
    x"00602825", -- 0x00001928
    x"8fc40040", -- 0x0000192c
    x"0c000565", -- 0x00001930
    x"00000000", -- 0x00001934
    x"02228821", -- 0x00001938
    x"10000062", -- 0x0000193c
    x"00000000", -- 0x00001940
    x"92030000", -- 0x00001944
    x"24020078", -- 0x00001948
    x"14620013", -- 0x0000194c
    x"00000000", -- 0x00001950
    x"8fc20044", -- 0x00001954
    x"00000000", -- 0x00001958
    x"24430004", -- 0x0000195c
    x"afc30044", -- 0x00001960
    x"8c430000", -- 0x00001964
    x"24020061", -- 0x00001968
    x"afa20018", -- 0x0000196c
    x"afb30014", -- 0x00001970
    x"afb20010", -- 0x00001974
    x"00003825", -- 0x00001978
    x"24060010", -- 0x0000197c
    x"00602825", -- 0x00001980
    x"8fc40040", -- 0x00001984
    x"0c000565", -- 0x00001988
    x"00000000", -- 0x0000198c
    x"02228821", -- 0x00001990
    x"1000004c", -- 0x00001994
    x"00000000", -- 0x00001998
    x"92030000", -- 0x0000199c
    x"24020058", -- 0x000019a0
    x"14620013", -- 0x000019a4
    x"00000000", -- 0x000019a8
    x"8fc20044", -- 0x000019ac
    x"00000000", -- 0x000019b0
    x"24430004", -- 0x000019b4
    x"afc30044", -- 0x000019b8
    x"8c430000", -- 0x000019bc
    x"24020041", -- 0x000019c0
    x"afa20018", -- 0x000019c4
    x"afb30014", -- 0x000019c8
    x"afb20010", -- 0x000019cc
    x"00003825", -- 0x000019d0
    x"24060010", -- 0x000019d4
    x"00602825", -- 0x000019d8
    x"8fc40040", -- 0x000019dc
    x"0c000565", -- 0x000019e0
    x"00000000", -- 0x000019e4
    x"02228821", -- 0x000019e8
    x"10000036", -- 0x000019ec
    x"00000000", -- 0x000019f0
    x"92030000", -- 0x000019f4
    x"24020075", -- 0x000019f8
    x"14620013", -- 0x000019fc
    x"00000000", -- 0x00001a00
    x"8fc20044", -- 0x00001a04
    x"00000000", -- 0x00001a08
    x"24430004", -- 0x00001a0c
    x"afc30044", -- 0x00001a10
    x"8c430000", -- 0x00001a14
    x"24020061", -- 0x00001a18
    x"afa20018", -- 0x00001a1c
    x"afb30014", -- 0x00001a20
    x"afb20010", -- 0x00001a24
    x"00003825", -- 0x00001a28
    x"2406000a", -- 0x00001a2c
    x"00602825", -- 0x00001a30
    x"8fc40040", -- 0x00001a34
    x"0c000565", -- 0x00001a38
    x"00000000", -- 0x00001a3c
    x"02228821", -- 0x00001a40
    x"10000020", -- 0x00001a44
    x"00000000", -- 0x00001a48
    x"92030000", -- 0x00001a4c
    x"24020063", -- 0x00001a50
    x"1462001c", -- 0x00001a54
    x"00000000", -- 0x00001a58
    x"8fc20044", -- 0x00001a5c
    x"00000000", -- 0x00001a60
    x"24430004", -- 0x00001a64
    x"afc30044", -- 0x00001a68
    x"8c420000", -- 0x00001a6c
    x"00000000", -- 0x00001a70
    x"304200ff", -- 0x00001a74
    x"a3c20020", -- 0x00001a78
    x"a3c00021", -- 0x00001a7c
    x"02603825", -- 0x00001a80
    x"02403025", -- 0x00001a84
    x"27c20020", -- 0x00001a88
    x"00402825", -- 0x00001a8c
    x"8fc40040", -- 0x00001a90
    x"0c0004f4", -- 0x00001a94
    x"00000000", -- 0x00001a98
    x"02228821", -- 0x00001a9c
    x"10000009", -- 0x00001aa0
    x"00000000", -- 0x00001aa4
    x"00000000", -- 0x00001aa8
    x"92020000", -- 0x00001aac
    x"00000000", -- 0x00001ab0
    x"00402825", -- 0x00001ab4
    x"8fc40040", -- 0x00001ab8
    x"0c0004cf", -- 0x00001abc
    x"00000000", -- 0x00001ac0
    x"26310001", -- 0x00001ac4
    x"26100001", -- 0x00001ac8
    x"92020000", -- 0x00001acc
    x"00000000", -- 0x00001ad0
    x"1440ff39", -- 0x00001ad4
    x"00000000", -- 0x00001ad8
    x"10000002", -- 0x00001adc
    x"00000000", -- 0x00001ae0
    x"00000000", -- 0x00001ae4
    x"8fc20040", -- 0x00001ae8
    x"00000000", -- 0x00001aec
    x"10400006", -- 0x00001af0
    x"00000000", -- 0x00001af4
    x"8fc20040", -- 0x00001af8
    x"00000000", -- 0x00001afc
    x"8c420000", -- 0x00001b00
    x"00000000", -- 0x00001b04
    x"a0400000", -- 0x00001b08
    x"02201025", -- 0x00001b0c
    x"03c0e825", -- 0x00001b10
    x"8fbf003c", -- 0x00001b14
    x"8fbe0038", -- 0x00001b18
    x"8fb30034", -- 0x00001b1c
    x"8fb20030", -- 0x00001b20
    x"8fb1002c", -- 0x00001b24
    x"8fb00028", -- 0x00001b28
    x"27bd0040", -- 0x00001b2c
    x"03e00008", -- 0x00001b30
    x"00000000", -- 0x00001b34
    x"27bdffe8", -- 0x00001b38
    x"afbf0014", -- 0x00001b3c
    x"afbe0010", -- 0x00001b40
    x"03a0f025", -- 0x00001b44
    x"afc40018", -- 0x00001b48
    x"afc5001c", -- 0x00001b4c
    x"afc60020", -- 0x00001b50
    x"afc70024", -- 0x00001b54
    x"27df0018", -- 0x00001b58
    x"03e02825", -- 0x00001b5c
    x"00002025", -- 0x00001b60
    x"0c0005db", -- 0x00001b64
    x"00000000", -- 0x00001b68
    x"03c0e825", -- 0x00001b6c
    x"8fbf0014", -- 0x00001b70
    x"8fbe0010", -- 0x00001b74
    x"27bd0018", -- 0x00001b78
    x"03e00008", -- 0x00001b7c
    x"00000000", -- 0x00001b80
    x"27bdffe8", -- 0x00001b84
    x"afbf0014", -- 0x00001b88
    x"afbe0010", -- 0x00001b8c
    x"03a0f025", -- 0x00001b90
    x"afc40018", -- 0x00001b94
    x"afc5001c", -- 0x00001b98
    x"afc60020", -- 0x00001b9c
    x"afc70024", -- 0x00001ba0
    x"27df001c", -- 0x00001ba4
    x"03e02825", -- 0x00001ba8
    x"27c40018", -- 0x00001bac
    x"0c0005db", -- 0x00001bb0
    x"00000000", -- 0x00001bb4
    x"03c0e825", -- 0x00001bb8
    x"8fbf0014", -- 0x00001bbc
    x"8fbe0010", -- 0x00001bc0
    x"27bd0018", -- 0x00001bc4
    x"03e00008", -- 0x00001bc8
    x"00000000", -- 0x00001bcc
    x"27bdfff8", -- 0x00001bd0
    x"afbe0004", -- 0x00001bd4
    x"03a0f025", -- 0x00001bd8
    x"afc40008", -- 0x00001bdc
    x"afc5000c", -- 0x00001be0
    x"afc60010", -- 0x00001be4
    x"afc70014", -- 0x00001be8
    x"8fc20008", -- 0x00001bec
    x"8fc3000c", -- 0x00001bf0
    x"00000000", -- 0x00001bf4
    x"ac430004", -- 0x00001bf8
    x"8fc20008", -- 0x00001bfc
    x"8fc30010", -- 0x00001c00
    x"00000000", -- 0x00001c04
    x"ac430008", -- 0x00001c08
    x"8fc20008", -- 0x00001c0c
    x"8fc30014", -- 0x00001c10
    x"00000000", -- 0x00001c14
    x"ac43000c", -- 0x00001c18
    x"8fc20008", -- 0x00001c1c
    x"8fc30018", -- 0x00001c20
    x"00000000", -- 0x00001c24
    x"ac430014", -- 0x00001c28
    x"00000000", -- 0x00001c2c
    x"03c0e825", -- 0x00001c30
    x"8fbe0004", -- 0x00001c34
    x"27bd0008", -- 0x00001c38
    x"03e00008", -- 0x00001c3c
    x"00000000", -- 0x00001c40
    x"27bdfff0", -- 0x00001c44
    x"afbe000c", -- 0x00001c48
    x"03a0f025", -- 0x00001c4c
    x"afc40010", -- 0x00001c50
    x"27820008", -- 0x00001c54
    x"afc20000", -- 0x00001c58
    x"1000000d", -- 0x00001c5c
    x"00000000", -- 0x00001c60
    x"8fc20000", -- 0x00001c64
    x"00000000", -- 0x00001c68
    x"8c430000", -- 0x00001c6c
    x"8fc20010", -- 0x00001c70
    x"00000000", -- 0x00001c74
    x"1062000e", -- 0x00001c78
    x"00000000", -- 0x00001c7c
    x"8fc20000", -- 0x00001c80
    x"00000000", -- 0x00001c84
    x"8c420000", -- 0x00001c88
    x"00000000", -- 0x00001c8c
    x"afc20000", -- 0x00001c90
    x"8fc20000", -- 0x00001c94
    x"00000000", -- 0x00001c98
    x"8c420000", -- 0x00001c9c
    x"00000000", -- 0x00001ca0
    x"1440ffef", -- 0x00001ca4
    x"00000000", -- 0x00001ca8
    x"10000002", -- 0x00001cac
    x"00000000", -- 0x00001cb0
    x"00000000", -- 0x00001cb4
    x"8fc20000", -- 0x00001cb8
    x"00000000", -- 0x00001cbc
    x"8c420000", -- 0x00001cc0
    x"00000000", -- 0x00001cc4
    x"1440000f", -- 0x00001cc8
    x"00000000", -- 0x00001ccc
    x"8fc20010", -- 0x00001cd0
    x"00000000", -- 0x00001cd4
    x"ac400000", -- 0x00001cd8
    x"8fc20010", -- 0x00001cdc
    x"00000000", -- 0x00001ce0
    x"8c43000c", -- 0x00001ce4
    x"8fc20010", -- 0x00001ce8
    x"00000000", -- 0x00001cec
    x"ac430010", -- 0x00001cf0
    x"8fc20000", -- 0x00001cf4
    x"8fc30010", -- 0x00001cf8
    x"00000000", -- 0x00001cfc
    x"ac430000", -- 0x00001d00
    x"00000000", -- 0x00001d04
    x"00000000", -- 0x00001d08
    x"03c0e825", -- 0x00001d0c
    x"8fbe000c", -- 0x00001d10
    x"27bd0010", -- 0x00001d14
    x"03e00008", -- 0x00001d18
    x"00000000", -- 0x00001d1c
    x"27bdfff0", -- 0x00001d20
    x"afbe000c", -- 0x00001d24
    x"03a0f025", -- 0x00001d28
    x"afc40010", -- 0x00001d2c
    x"afc00004", -- 0x00001d30
    x"27820008", -- 0x00001d34
    x"afc20000", -- 0x00001d38
    x"10000019", -- 0x00001d3c
    x"00000000", -- 0x00001d40
    x"8fc20000", -- 0x00001d44
    x"00000000", -- 0x00001d48
    x"8c430000", -- 0x00001d4c
    x"8fc20010", -- 0x00001d50
    x"00000000", -- 0x00001d54
    x"1462000d", -- 0x00001d58
    x"00000000", -- 0x00001d5c
    x"8fc20000", -- 0x00001d60
    x"00000000", -- 0x00001d64
    x"8c420000", -- 0x00001d68
    x"00000000", -- 0x00001d6c
    x"8c430000", -- 0x00001d70
    x"8fc20000", -- 0x00001d74
    x"00000000", -- 0x00001d78
    x"ac430000", -- 0x00001d7c
    x"24020001", -- 0x00001d80
    x"afc20004", -- 0x00001d84
    x"1000000c", -- 0x00001d88
    x"00000000", -- 0x00001d8c
    x"8fc20000", -- 0x00001d90
    x"00000000", -- 0x00001d94
    x"8c420000", -- 0x00001d98
    x"00000000", -- 0x00001d9c
    x"afc20000", -- 0x00001da0
    x"8fc20000", -- 0x00001da4
    x"00000000", -- 0x00001da8
    x"8c420000", -- 0x00001dac
    x"00000000", -- 0x00001db0
    x"1440ffe3", -- 0x00001db4
    x"00000000", -- 0x00001db8
    x"8fc20004", -- 0x00001dbc
    x"03c0e825", -- 0x00001dc0
    x"8fbe000c", -- 0x00001dc4
    x"27bd0010", -- 0x00001dc8
    x"03e00008", -- 0x00001dcc
    x"00000000", -- 0x00001dd0
    x"27bdffe0", -- 0x00001dd4
    x"afbf001c", -- 0x00001dd8
    x"afbe0018", -- 0x00001ddc
    x"03a0f025", -- 0x00001de0
    x"afc40020", -- 0x00001de4
    x"8f830090", -- 0x00001de8
    x"8fc20020", -- 0x00001dec
    x"00000000", -- 0x00001df0
    x"00621021", -- 0x00001df4
    x"af820090", -- 0x00001df8
    x"8f820090", -- 0x00001dfc
    x"00000000", -- 0x00001e00
    x"24420001", -- 0x00001e04
    x"af820090", -- 0x00001e08
    x"8fc30020", -- 0x00001e0c
    x"00000000", -- 0x00001e10
    x"0043102b", -- 0x00001e14
    x"10400005", -- 0x00001e18
    x"00000000", -- 0x00001e1c
    x"8f820094", -- 0x00001e20
    x"00000000", -- 0x00001e24
    x"24420001", -- 0x00001e28
    x"af820094", -- 0x00001e2c
    x"27820008", -- 0x00001e30
    x"afc20010", -- 0x00001e34
    x"10000056", -- 0x00001e38
    x"00000000", -- 0x00001e3c
    x"8fc20010", -- 0x00001e40
    x"00000000", -- 0x00001e44
    x"8c420000", -- 0x00001e48
    x"8fc30010", -- 0x00001e4c
    x"00000000", -- 0x00001e50
    x"8c630000", -- 0x00001e54
    x"00000000", -- 0x00001e58
    x"8c630010", -- 0x00001e5c
    x"00000000", -- 0x00001e60
    x"00602025", -- 0x00001e64
    x"8fc30020", -- 0x00001e68
    x"00000000", -- 0x00001e6c
    x"00831823", -- 0x00001e70
    x"ac430010", -- 0x00001e74
    x"8fc20010", -- 0x00001e78
    x"00000000", -- 0x00001e7c
    x"8c420000", -- 0x00001e80
    x"00000000", -- 0x00001e84
    x"8c420010", -- 0x00001e88
    x"00000000", -- 0x00001e8c
    x"1c400032", -- 0x00001e90
    x"00000000", -- 0x00001e94
    x"8fc20010", -- 0x00001e98
    x"00000000", -- 0x00001e9c
    x"8c420000", -- 0x00001ea0
    x"00000000", -- 0x00001ea4
    x"8c420004", -- 0x00001ea8
    x"8fc30010", -- 0x00001eac
    x"00000000", -- 0x00001eb0
    x"8c630000", -- 0x00001eb4
    x"00000000", -- 0x00001eb8
    x"8c630008", -- 0x00001ebc
    x"00000000", -- 0x00001ec0
    x"00602025", -- 0x00001ec4
    x"0040f809", -- 0x00001ec8
    x"00000000", -- 0x00001ecc
    x"8fc20010", -- 0x00001ed0
    x"00000000", -- 0x00001ed4
    x"8c420000", -- 0x00001ed8
    x"00000000", -- 0x00001edc
    x"8c420014", -- 0x00001ee0
    x"24030001", -- 0x00001ee4
    x"1043000e", -- 0x00001ee8
    x"00000000", -- 0x00001eec
    x"24030002", -- 0x00001ef0
    x"14430019", -- 0x00001ef4
    x"00000000", -- 0x00001ef8
    x"8fc20010", -- 0x00001efc
    x"00000000", -- 0x00001f00
    x"8c420000", -- 0x00001f04
    x"00000000", -- 0x00001f08
    x"8c430000", -- 0x00001f0c
    x"8fc20010", -- 0x00001f10
    x"00000000", -- 0x00001f14
    x"ac430000", -- 0x00001f18
    x"1000000f", -- 0x00001f1c
    x"00000000", -- 0x00001f20
    x"8fc20010", -- 0x00001f24
    x"00000000", -- 0x00001f28
    x"8c420000", -- 0x00001f2c
    x"00000000", -- 0x00001f30
    x"8c43000c", -- 0x00001f34
    x"8fc20010", -- 0x00001f38
    x"00000000", -- 0x00001f3c
    x"8c420000", -- 0x00001f40
    x"00000000", -- 0x00001f44
    x"8c440010", -- 0x00001f48
    x"00000000", -- 0x00001f4c
    x"00831821", -- 0x00001f50
    x"ac430010", -- 0x00001f54
    x"00000000", -- 0x00001f58
    x"8fc20010", -- 0x00001f5c
    x"00000000", -- 0x00001f60
    x"8c420000", -- 0x00001f64
    x"00000000", -- 0x00001f68
    x"10400006", -- 0x00001f6c
    x"00000000", -- 0x00001f70
    x"8fc20010", -- 0x00001f74
    x"00000000", -- 0x00001f78
    x"8c420000", -- 0x00001f7c
    x"10000003", -- 0x00001f80
    x"00000000", -- 0x00001f84
    x"8fc20010", -- 0x00001f88
    x"00000000", -- 0x00001f8c
    x"afc20010", -- 0x00001f90
    x"8fc20010", -- 0x00001f94
    x"00000000", -- 0x00001f98
    x"8c420000", -- 0x00001f9c
    x"00000000", -- 0x00001fa0
    x"1440ffa6", -- 0x00001fa4
    x"00000000", -- 0x00001fa8
    x"00000000", -- 0x00001fac
    x"03c0e825", -- 0x00001fb0
    x"8fbf001c", -- 0x00001fb4
    x"8fbe0018", -- 0x00001fb8
    x"27bd0020", -- 0x00001fbc
    x"03e00008", -- 0x00001fc0
    x"00000000", -- 0x00001fc4
    x"27bdfff0", -- 0x00001fc8
    x"afbe000c", -- 0x00001fcc
    x"03a0f025", -- 0x00001fd0
    x"afc40010", -- 0x00001fd4
    x"8fc20010", -- 0x00001fd8
    x"00000000", -- 0x00001fdc
    x"1040000f", -- 0x00001fe0
    x"00000000", -- 0x00001fe4
    x"8f830090", -- 0x00001fe8
    x"8fc20010", -- 0x00001fec
    x"00000000", -- 0x00001ff0
    x"00621021", -- 0x00001ff4
    x"afc20000", -- 0x00001ff8
    x"00000000", -- 0x00001ffc
    x"8f830090", -- 0x00002000
    x"8fc20000", -- 0x00002004
    x"00000000", -- 0x00002008
    x"1462fffc", -- 0x0000200c
    x"00000000", -- 0x00002010
    x"00000000", -- 0x00002014
    x"10000002", -- 0x00002018
    x"00000000", -- 0x0000201c
    x"00000000", -- 0x00002020
    x"03c0e825", -- 0x00002024
    x"8fbe000c", -- 0x00002028
    x"27bd0010", -- 0x0000202c
    x"03e00008", -- 0x00002030
    x"00000000", -- 0x00002034
    x"27bdffe8", -- 0x00002038
    x"afbf0014", -- 0x0000203c
    x"afbe0010", -- 0x00002040
    x"03a0f025", -- 0x00002044
    x"afc40018", -- 0x00002048
    x"afc5001c", -- 0x0000204c
    x"afc60020", -- 0x00002050
    x"afc70024", -- 0x00002054
    x"8fc20018", -- 0x00002058
    x"00000000", -- 0x0000205c
    x"af82000c", -- 0x00002060
    x"8f82000c", -- 0x00002064
    x"00000000", -- 0x00002068
    x"24460008", -- 0x0000206c
    x"8fc20028", -- 0x00002070
    x"00000000", -- 0x00002074
    x"00021d80", -- 0x00002078
    x"8fc20024", -- 0x0000207c
    x"00000000", -- 0x00002080
    x"00021500", -- 0x00002084
    x"00621825", -- 0x00002088
    x"8fc20020", -- 0x0000208c
    x"00000000", -- 0x00002090
    x"2442ffff", -- 0x00002094
    x"00021400", -- 0x00002098
    x"00621825", -- 0x0000209c
    x"3c0202fa", -- 0x000020a0
    x"3444f080", -- 0x000020a4
    x"8fc2001c", -- 0x000020a8
    x"00000000", -- 0x000020ac
    x"0082001b", -- 0x000020b0
    x"00001010", -- 0x000020b4
    x"00001012", -- 0x000020b8
    x"2442ffff", -- 0x000020bc
    x"00621825", -- 0x000020c0
    x"3c020100", -- 0x000020c4
    x"00621025", -- 0x000020c8
    x"00402825", -- 0x000020cc
    x"00c02025", -- 0x000020d0
    x"0c00012b", -- 0x000020d4
    x"00000000", -- 0x000020d8
    x"00000000", -- 0x000020dc
    x"03c0e825", -- 0x000020e0
    x"8fbf0014", -- 0x000020e4
    x"8fbe0010", -- 0x000020e8
    x"27bd0018", -- 0x000020ec
    x"03e00008", -- 0x000020f0
    x"00000000", -- 0x000020f4
    x"27bdffe0", -- 0x000020f8
    x"afbf001c", -- 0x000020fc
    x"afbe0018", -- 0x00002100
    x"03a0f025", -- 0x00002104
    x"27c20010", -- 0x00002108
    x"00402825", -- 0x0000210c
    x"3c020000", -- 0x00002110
    x"24444010", -- 0x00002114
    x"0c0000d5", -- 0x00002118
    x"00000000", -- 0x0000211c
    x"00401825", -- 0x00002120
    x"2402ffff", -- 0x00002124
    x"14620004", -- 0x00002128
    x"00000000", -- 0x0000212c
    x"2402ffff", -- 0x00002130
    x"10000002", -- 0x00002134
    x"00000000", -- 0x00002138
    x"93c20010", -- 0x0000213c
    x"03c0e825", -- 0x00002140
    x"8fbf001c", -- 0x00002144
    x"8fbe0018", -- 0x00002148
    x"27bd0020", -- 0x0000214c
    x"03e00008", -- 0x00002150
    x"00000000", -- 0x00002154
    x"27bdffe0", -- 0x00002158
    x"afbf001c", -- 0x0000215c
    x"afbe0018", -- 0x00002160
    x"afb00014", -- 0x00002164
    x"03a0f025", -- 0x00002168
    x"afc40020", -- 0x0000216c
    x"8fc50020", -- 0x00002170
    x"3c020000", -- 0x00002174
    x"24444070", -- 0x00002178
    x"0c00007e", -- 0x0000217c
    x"00000000", -- 0x00002180
    x"8f82000c", -- 0x00002184
    x"00000000", -- 0x00002188
    x"24500008", -- 0x0000218c
    x"8f82000c", -- 0x00002190
    x"00000000", -- 0x00002194
    x"24420008", -- 0x00002198
    x"00402025", -- 0x0000219c
    x"0c00013a", -- 0x000021a0
    x"00000000", -- 0x000021a4
    x"00401825", -- 0x000021a8
    x"3c020200", -- 0x000021ac
    x"00621025", -- 0x000021b0
    x"00402825", -- 0x000021b4
    x"02002025", -- 0x000021b8
    x"0c00012b", -- 0x000021bc
    x"00000000", -- 0x000021c0
    x"00000000", -- 0x000021c4
    x"03c0e825", -- 0x000021c8
    x"8fbf001c", -- 0x000021cc
    x"8fbe0018", -- 0x000021d0
    x"8fb00014", -- 0x000021d4
    x"27bd0020", -- 0x000021d8
    x"03e00008", -- 0x000021dc
    x"00000000", -- 0x000021e0
    x"00000000", -- 0x000021e4
    x"02200000", -- 0x000021e8
    x"01000101", -- 0x000021ec
    x"00000000", -- 0x000021f0
    x"00000000", -- 0x000021f4
    x"00000001", -- 0x000021f8
    x"00000000", -- 0x000021fc
    x"6c756e28", -- 0x00002200
    x"0000296c", -- 0x00002204
    x"00000000", -- 0x00002208
    x"00000000", -- 0x0000220c
    x"00000000", -- 0x00002210
    x"00000000", -- 0x00002214
    x"00000000", -- 0x00002218
    x"00000000", -- 0x0000221c
    x"00000000", -- 0x00002220
    x"00000000", -- 0x00002224
    x"00000000", -- 0x00002228
    x"00000000", -- 0x0000222c
    x"00000000", -- 0x00002230
    x"00000000", -- 0x00002234
    x"00000000", -- 0x00002238
    x"00000000", -- 0x0000223c
    x"00000000", -- 0x00002240
    x"00000000", -- 0x00002244
    x"00000000", -- 0x00002248
    x"00000000", -- 0x0000224c
    x"00000000", -- 0x00002250
    x"00000000", -- 0x00002254
    x"00000000", -- 0x00002258
    x"00000000", -- 0x0000225c
    x"00000000", -- 0x00002260
    x"00000000", -- 0x00002264
    x"00000000", -- 0x00002268
    x"00000000", -- 0x0000226c
    x"00000000", -- 0x00002270
    x"00000000", -- 0x00002274
    x"00000000", -- 0x00002278
    x"00000000", -- 0x0000227c
    x"00000000", -- 0x00002280
    x"00000000", -- 0x00002284
    x"00000000", -- 0x00002288
    x"00000000", -- 0x0000228c
    x"00000000", -- 0x00002290
    x"00000000", -- 0x00002294
    x"00000000", -- 0x00002298
    x"00000000", -- 0x0000229c
    x"00000000", -- 0x000022a0
    x"00000000", -- 0x000022a4
    x"00000000", -- 0x000022a8
    x"00000000", -- 0x000022ac
    x"00000000", -- 0x000022b0
    x"00000000", -- 0x000022b4
    x"00000000", -- 0x000022b8
    x"00000000", -- 0x000022bc
    x"00000000", -- 0x000022c0
    x"00000000", -- 0x000022c4
    x"00000000", -- 0x000022c8
    x"00000000", -- 0x000022cc
    x"00000000", -- 0x000022d0
    x"00000000", -- 0x000022d4
    x"00000000", -- 0x000022d8
    x"00000000", -- 0x000022dc
    x"00000000", -- 0x000022e0
    x"00000000", -- 0x000022e4
    x"00000000", -- 0x000022e8
    x"00000000", -- 0x000022ec
    x"00000000", -- 0x000022f0
    x"00000000", -- 0x000022f4
    x"00000000", -- 0x000022f8
    x"00000000", -- 0x000022fc
    x"00000000", -- 0x00002300
    x"00000000", -- 0x00002304
    x"00000000", -- 0x00002308
    x"00000000", -- 0x0000230c
    x"00000000", -- 0x00002310
    x"00000000", -- 0x00002314
    x"00000000", -- 0x00002318
    x"00000000", -- 0x0000231c
    x"00000000", -- 0x00002320
    x"00000000", -- 0x00002324
    x"00000000", -- 0x00002328
    x"00000000", -- 0x0000232c
    x"00000000", -- 0x00002330
    x"00000000", -- 0x00002334
    x"00000000", -- 0x00002338
    x"00000000", -- 0x0000233c
    x"00000000", -- 0x00002340
    x"00000000", -- 0x00002344
    x"00000000", -- 0x00002348
    x"00000000", -- 0x0000234c
    x"00000000", -- 0x00002350
    x"00000000", -- 0x00002354
    x"00000000", -- 0x00002358
    x"00000000", -- 0x0000235c
    x"00000000", -- 0x00002360
    x"00000000", -- 0x00002364
    x"00000000", -- 0x00002368
    x"00000000", -- 0x0000236c
    x"00000000", -- 0x00002370
    x"00000000", -- 0x00002374
    x"00000000", -- 0x00002378
    x"00000000", -- 0x0000237c
    x"00000000", -- 0x00002380
    x"00000000", -- 0x00002384
    x"00000000", -- 0x00002388
    x"00000000", -- 0x0000238c
    x"00000000", -- 0x00002390
    x"00000000", -- 0x00002394
    x"00000000", -- 0x00002398
    x"00000000", -- 0x0000239c
    x"00000000", -- 0x000023a0
    x"00000000", -- 0x000023a4
    x"00000000", -- 0x000023a8
    x"00000000", -- 0x000023ac
    x"00000000", -- 0x000023b0
    x"00000000", -- 0x000023b4
    x"00000000", -- 0x000023b8
    x"00000000", -- 0x000023bc
    x"00000000", -- 0x000023c0
    x"00000000", -- 0x000023c4
    x"00000000", -- 0x000023c8
    x"00000000", -- 0x000023cc
    x"00000000", -- 0x000023d0
    x"00000000", -- 0x000023d4
    x"00000000", -- 0x000023d8
    x"00000000", -- 0x000023dc
    x"00000000", -- 0x000023e0
    x"00000000", -- 0x000023e4
    x"00000000", -- 0x000023e8
    x"00000000", -- 0x000023ec
    x"00000000", -- 0x000023f0
    x"00000000", -- 0x000023f4
    x"00000000", -- 0x000023f8
    x"00000000", -- 0x000023fc
    x"00000000", -- 0x00002400
    x"00000000", -- 0x00002404
    x"00000000", -- 0x00002408
    x"00000000", -- 0x0000240c
    x"00000000", -- 0x00002410
    x"00000000", -- 0x00002414
    x"00000000", -- 0x00002418
    x"00000000", -- 0x0000241c
    x"00000000", -- 0x00002420
    x"00000000", -- 0x00002424
    x"00000000", -- 0x00002428
    x"00000000", -- 0x0000242c
    x"00000000", -- 0x00002430
    x"00000000", -- 0x00002434
    x"00000000", -- 0x00002438
    x"00000000", -- 0x0000243c
    x"00000000", -- 0x00002440
    x"00000000", -- 0x00002444
    x"00000000", -- 0x00002448
    x"00000000", -- 0x0000244c
    x"00000000", -- 0x00002450
    x"00000000", -- 0x00002454
    x"00000000", -- 0x00002458
    x"00000000", -- 0x0000245c
    x"00000000", -- 0x00002460
    x"00000000", -- 0x00002464
    x"00000000", -- 0x00002468
    x"00000000", -- 0x0000246c
    x"00000000", -- 0x00002470
    x"00000000", -- 0x00002474
    x"00000000", -- 0x00002478
    x"00000000", -- 0x0000247c
    x"00000000", -- 0x00002480
    x"00000000", -- 0x00002484
    x"00000000", -- 0x00002488
    x"00000000", -- 0x0000248c
    x"00000000", -- 0x00002490
    x"00000000", -- 0x00002494
    x"00000000", -- 0x00002498
    x"00000000", -- 0x0000249c
    x"00000000", -- 0x000024a0
    x"00000000", -- 0x000024a4
    x"00000000", -- 0x000024a8
    x"00000000", -- 0x000024ac
    x"00000000", -- 0x000024b0
    x"00000000", -- 0x000024b4
    x"00000000", -- 0x000024b8
    x"00000000", -- 0x000024bc
    x"00000000", -- 0x000024c0
    x"00000000", -- 0x000024c4
    x"00000000", -- 0x000024c8
    x"00000000", -- 0x000024cc
    x"00000000", -- 0x000024d0
    x"00000000", -- 0x000024d4
    x"00000000", -- 0x000024d8
    x"00000000", -- 0x000024dc
    x"00000000", -- 0x000024e0
    x"00000000", -- 0x000024e4
    x"00000000", -- 0x000024e8
    x"00000000", -- 0x000024ec
    x"00000000", -- 0x000024f0
    x"00000000", -- 0x000024f4
    x"00000000", -- 0x000024f8
    x"00000000", -- 0x000024fc
    x"00000000", -- 0x00002500
    x"00000000", -- 0x00002504
    x"00000000", -- 0x00002508
    x"00000000", -- 0x0000250c
    x"00000000", -- 0x00002510
    x"00000000", -- 0x00002514
    x"00000000", -- 0x00002518
    x"00000000", -- 0x0000251c
    x"00000000", -- 0x00002520
    x"00000000", -- 0x00002524
    x"00000000", -- 0x00002528
    x"00000000", -- 0x0000252c
    x"00000000", -- 0x00002530
    x"00000000", -- 0x00002534
    x"00000000", -- 0x00002538
    x"00000000", -- 0x0000253c
    x"00000000", -- 0x00002540
    x"00000000", -- 0x00002544
    x"00000000", -- 0x00002548
    x"00000000", -- 0x0000254c
    x"00000000", -- 0x00002550
    x"00000000", -- 0x00002554
    x"00000000", -- 0x00002558
    x"00000000", -- 0x0000255c
    x"00000000", -- 0x00002560
    x"00000000", -- 0x00002564
    x"00000000", -- 0x00002568
    x"00000000", -- 0x0000256c
    x"00000000", -- 0x00002570
    x"00000000", -- 0x00002574
    x"00000000", -- 0x00002578
    x"00000000", -- 0x0000257c
    x"00000000", -- 0x00002580
    x"00000000", -- 0x00002584
    x"00000000", -- 0x00002588
    x"00000000", -- 0x0000258c
    x"00000000", -- 0x00002590
    x"00000000", -- 0x00002594
    x"00000000", -- 0x00002598
    x"00000000", -- 0x0000259c
    x"00000000", -- 0x000025a0
    x"00000000", -- 0x000025a4
    x"00000000", -- 0x000025a8
    x"00000000", -- 0x000025ac
    x"00000000", -- 0x000025b0
    x"00000000", -- 0x000025b4
    x"00000000", -- 0x000025b8
    x"00000000", -- 0x000025bc
    x"00000000", -- 0x000025c0
    x"00000000", -- 0x000025c4
    x"00000000", -- 0x000025c8
    x"00000000", -- 0x000025cc
    x"00000000", -- 0x000025d0
    x"00000000", -- 0x000025d4
    x"00000000", -- 0x000025d8
    x"00000000", -- 0x000025dc
    x"00000000", -- 0x000025e0
    x"00000000", -- 0x000025e4
    x"00000000", -- 0x000025e8
    x"00000000", -- 0x000025ec
    x"00000000", -- 0x000025f0
    x"00000000", -- 0x000025f4
    x"00000000", -- 0x000025f8
    x"00000000", -- 0x000025fc
    x"00000000", -- 0x00002600
    x"00000000", -- 0x00002604
    x"00000000", -- 0x00002608
    x"00000000", -- 0x0000260c
    x"00000000", -- 0x00002610
    x"00000000", -- 0x00002614
    x"00000000", -- 0x00002618
    x"00000000", -- 0x0000261c
    x"00000000", -- 0x00002620
    x"00000000", -- 0x00002624
    x"00000000", -- 0x00002628
    x"00000000", -- 0x0000262c
    x"00000000", -- 0x00002630
    x"00000000", -- 0x00002634
    x"00000000", -- 0x00002638
    x"00000000", -- 0x0000263c
    x"00000000", -- 0x00002640
    x"00000000", -- 0x00002644
    x"00000000", -- 0x00002648
    x"00000000", -- 0x0000264c
    x"00000000", -- 0x00002650
    x"00000000", -- 0x00002654
    x"00000000", -- 0x00002658
    x"00000000", -- 0x0000265c
    x"00000000", -- 0x00002660
    x"00000000", -- 0x00002664
    x"00000000", -- 0x00002668
    x"00000000", -- 0x0000266c
    x"00000000", -- 0x00002670
    x"00000000", -- 0x00002674
    x"00000000", -- 0x00002678
    x"00000000", -- 0x0000267c
    x"00000000", -- 0x00002680
    x"00000000", -- 0x00002684
    x"00000000", -- 0x00002688
    x"00000000", -- 0x0000268c
    x"00000000", -- 0x00002690
    x"00000000", -- 0x00002694
    x"00000000", -- 0x00002698
    x"00000000", -- 0x0000269c
    x"00000000", -- 0x000026a0
    x"00000000", -- 0x000026a4
    x"00000000", -- 0x000026a8
    x"00000000", -- 0x000026ac
    x"00000000", -- 0x000026b0
    x"00000000", -- 0x000026b4
    x"00000000", -- 0x000026b8
    x"00000000", -- 0x000026bc
    x"00000000", -- 0x000026c0
    x"00000000", -- 0x000026c4
    x"00000000", -- 0x000026c8
    x"00000000", -- 0x000026cc
    x"00000000", -- 0x000026d0
    x"00000000", -- 0x000026d4
    x"00000000", -- 0x000026d8
    x"00000000", -- 0x000026dc
    x"00000000", -- 0x000026e0
    x"00000000", -- 0x000026e4
    x"00000000", -- 0x000026e8
    x"00000000", -- 0x000026ec
    x"00000000", -- 0x000026f0
    x"00000000", -- 0x000026f4
    x"00000000", -- 0x000026f8
    x"00000000", -- 0x000026fc
    x"00000000", -- 0x00002700
    x"00000000", -- 0x00002704
    x"00000000", -- 0x00002708
    x"00000000", -- 0x0000270c
    x"00000000", -- 0x00002710
    x"00000000", -- 0x00002714
    x"00000000", -- 0x00002718
    x"00000000", -- 0x0000271c
    x"00000000", -- 0x00002720
    x"00000000", -- 0x00002724
    x"00000000", -- 0x00002728
    x"00000000", -- 0x0000272c
    x"00000000", -- 0x00002730
    x"00000000", -- 0x00002734
    x"00000000", -- 0x00002738
    x"00000000", -- 0x0000273c
    x"00000000", -- 0x00002740
    x"00000000", -- 0x00002744
    x"00000000", -- 0x00002748
    x"00000000", -- 0x0000274c
    x"00000000", -- 0x00002750
    x"00000000", -- 0x00002754
    x"00000000", -- 0x00002758
    x"00000000", -- 0x0000275c
    x"00000000", -- 0x00002760
    x"00000000", -- 0x00002764
    x"00000000", -- 0x00002768
    x"00000000", -- 0x0000276c
    x"00000000", -- 0x00002770
    x"00000000", -- 0x00002774
    x"00000000", -- 0x00002778
    x"00000000", -- 0x0000277c
    x"00000000", -- 0x00002780
    x"00000000", -- 0x00002784
    x"00000000", -- 0x00002788
    x"00000000", -- 0x0000278c
    x"00000000", -- 0x00002790
    x"00000000", -- 0x00002794
    x"00000000", -- 0x00002798
    x"00000000", -- 0x0000279c
    x"00000000", -- 0x000027a0
    x"00000000", -- 0x000027a4
    x"00000000", -- 0x000027a8
    x"00000000", -- 0x000027ac
    x"00000000", -- 0x000027b0
    x"00000000", -- 0x000027b4
    x"00000000", -- 0x000027b8
    x"00000000", -- 0x000027bc
    x"00000000", -- 0x000027c0
    x"00000000", -- 0x000027c4
    x"00000000", -- 0x000027c8
    x"00000000", -- 0x000027cc
    x"00000000", -- 0x000027d0
    x"00000000", -- 0x000027d4
    x"00000000", -- 0x000027d8
    x"00000000", -- 0x000027dc
    x"00000000", -- 0x000027e0
    x"00000000", -- 0x000027e4
    x"00000000", -- 0x000027e8
    x"00000000", -- 0x000027ec
    x"00000000", -- 0x000027f0
    x"00000000", -- 0x000027f4
    x"00000000", -- 0x000027f8
    x"00000000", -- 0x000027fc
    x"00000000", -- 0x00002800
    x"00000000", -- 0x00002804
    x"00000000", -- 0x00002808
    x"00000000", -- 0x0000280c
    x"00000000", -- 0x00002810
    x"00000000", -- 0x00002814
    x"00000000", -- 0x00002818
    x"00000000", -- 0x0000281c
    x"00000000", -- 0x00002820
    x"00000000", -- 0x00002824
    x"00000000", -- 0x00002828
    x"00000000", -- 0x0000282c
    x"00000000", -- 0x00002830
    x"00000000", -- 0x00002834
    x"00000000", -- 0x00002838
    x"00000000", -- 0x0000283c
    x"00000000", -- 0x00002840
    x"00000000", -- 0x00002844
    x"00000000", -- 0x00002848
    x"00000000", -- 0x0000284c
    x"00000000", -- 0x00002850
    x"00000000", -- 0x00002854
    x"00000000", -- 0x00002858
    x"00000000", -- 0x0000285c
    x"00000000", -- 0x00002860
    x"00000000", -- 0x00002864
    x"00000000", -- 0x00002868
    x"00000000", -- 0x0000286c
    x"00000000", -- 0x00002870
    x"00000000", -- 0x00002874
    x"00000000", -- 0x00002878
    x"00000000", -- 0x0000287c
    x"00000000", -- 0x00002880
    x"00000000", -- 0x00002884
    x"00000000", -- 0x00002888
    x"00000000", -- 0x0000288c
    x"00000000", -- 0x00002890
    x"00000000", -- 0x00002894
    x"00000000", -- 0x00002898
    x"00000000", -- 0x0000289c
    x"00000000", -- 0x000028a0
    x"00000000", -- 0x000028a4
    x"00000000", -- 0x000028a8
    x"00000000", -- 0x000028ac
    x"00000000", -- 0x000028b0
    x"00000000", -- 0x000028b4
    x"00000000", -- 0x000028b8
    x"00000000", -- 0x000028bc
    x"00000000", -- 0x000028c0
    x"00000000", -- 0x000028c4
    x"00000000", -- 0x000028c8
    x"00000000", -- 0x000028cc
    x"00000000", -- 0x000028d0
    x"00000000", -- 0x000028d4
    x"00000000", -- 0x000028d8
    x"00000000", -- 0x000028dc
    x"00000000", -- 0x000028e0
    x"00000000", -- 0x000028e4
    x"00000000", -- 0x000028e8
    x"00000000", -- 0x000028ec
    x"00000000", -- 0x000028f0
    x"00000000", -- 0x000028f4
    x"00000000", -- 0x000028f8
    x"00000000", -- 0x000028fc
    x"00000000", -- 0x00002900
    x"00000000", -- 0x00002904
    x"00000000", -- 0x00002908
    x"00000000", -- 0x0000290c
    x"00000000", -- 0x00002910
    x"00000000", -- 0x00002914
    x"00000000", -- 0x00002918
    x"00000000", -- 0x0000291c
    x"00000000", -- 0x00002920
    x"00000000", -- 0x00002924
    x"00000000", -- 0x00002928
    x"00000000", -- 0x0000292c
    x"00000000", -- 0x00002930
    x"00000000", -- 0x00002934
    x"00000000", -- 0x00002938
    x"00000000", -- 0x0000293c
    x"00000000", -- 0x00002940
    x"00000000", -- 0x00002944
    x"00000000", -- 0x00002948
    x"00000000", -- 0x0000294c
    x"00000000", -- 0x00002950
    x"00000000", -- 0x00002954
    x"00000000", -- 0x00002958
    x"00000000", -- 0x0000295c
    x"00000000", -- 0x00002960
    x"00000000", -- 0x00002964
    x"00000000", -- 0x00002968
    x"00000000", -- 0x0000296c
    x"00000000", -- 0x00002970
    x"00000000", -- 0x00002974
    x"00000000", -- 0x00002978
    x"00000000", -- 0x0000297c
    x"00000000", -- 0x00002980
    x"00000000", -- 0x00002984
    x"00000000", -- 0x00002988
    x"00000000", -- 0x0000298c
    x"00000000", -- 0x00002990
    x"00000000", -- 0x00002994
    x"00000000", -- 0x00002998
    x"00000000", -- 0x0000299c
    x"00000000", -- 0x000029a0
    x"00000000", -- 0x000029a4
    x"00000000", -- 0x000029a8
    x"00000000", -- 0x000029ac
    x"00000000", -- 0x000029b0
    x"00000000", -- 0x000029b4
    x"00000000", -- 0x000029b8
    x"00000000", -- 0x000029bc
    x"00000000", -- 0x000029c0
    x"00000000", -- 0x000029c4
    x"00000000", -- 0x000029c8
    x"00000000", -- 0x000029cc
    x"00000000", -- 0x000029d0
    x"00000000", -- 0x000029d4
    x"00000000", -- 0x000029d8
    x"00000000", -- 0x000029dc
    x"00000000", -- 0x000029e0
    x"00000000", -- 0x000029e4
    x"00000000", -- 0x000029e8
    x"00000000", -- 0x000029ec
    x"00000000", -- 0x000029f0
    x"00000000", -- 0x000029f4
    x"00000000", -- 0x000029f8
    x"00000000", -- 0x000029fc
    x"00000000", -- 0x00002a00
    x"00000000", -- 0x00002a04
    x"00000000", -- 0x00002a08
    x"00000000", -- 0x00002a0c
    x"00000000", -- 0x00002a10
    x"00000000", -- 0x00002a14
    x"00000000", -- 0x00002a18
    x"00000000", -- 0x00002a1c
    x"00000000", -- 0x00002a20
    x"00000000", -- 0x00002a24
    x"00000000", -- 0x00002a28
    x"00000000", -- 0x00002a2c
    x"00000000", -- 0x00002a30
    x"00000000", -- 0x00002a34
    x"00000000", -- 0x00002a38
    x"00000000", -- 0x00002a3c
    x"00000000", -- 0x00002a40
    x"00000000", -- 0x00002a44
    x"00000000", -- 0x00002a48
    x"00000000", -- 0x00002a4c
    x"00000000", -- 0x00002a50
    x"00000000", -- 0x00002a54
    x"00000000", -- 0x00002a58
    x"00000000", -- 0x00002a5c
    x"00000000", -- 0x00002a60
    x"00000000", -- 0x00002a64
    x"00000000", -- 0x00002a68
    x"00000000", -- 0x00002a6c
    x"00000000", -- 0x00002a70
    x"00000000", -- 0x00002a74
    x"00000000", -- 0x00002a78
    x"00000000", -- 0x00002a7c
    x"00000000", -- 0x00002a80
    x"00000000", -- 0x00002a84
    x"00000000", -- 0x00002a88
    x"00000000", -- 0x00002a8c
    x"00000000", -- 0x00002a90
    x"00000000", -- 0x00002a94
    x"00000000", -- 0x00002a98
    x"00000000", -- 0x00002a9c
    x"00000000", -- 0x00002aa0
    x"00000000", -- 0x00002aa4
    x"00000000", -- 0x00002aa8
    x"00000000", -- 0x00002aac
    x"00000000", -- 0x00002ab0
    x"00000000", -- 0x00002ab4
    x"00000000", -- 0x00002ab8
    x"00000000", -- 0x00002abc
    x"00000000", -- 0x00002ac0
    x"00000000", -- 0x00002ac4
    x"00000000", -- 0x00002ac8
    x"00000000", -- 0x00002acc
    x"00000000", -- 0x00002ad0
    x"00000000", -- 0x00002ad4
    x"00000000", -- 0x00002ad8
    x"00000000", -- 0x00002adc
    x"00000000", -- 0x00002ae0
    x"00000000", -- 0x00002ae4
    x"00000000", -- 0x00002ae8
    x"00000000", -- 0x00002aec
    x"00000000", -- 0x00002af0
    x"00000000", -- 0x00002af4
    x"00000000", -- 0x00002af8
    x"00000000", -- 0x00002afc
    x"00000000", -- 0x00002b00
    x"00000000", -- 0x00002b04
    x"00000000", -- 0x00002b08
    x"00000000", -- 0x00002b0c
    x"00000000", -- 0x00002b10
    x"00000000", -- 0x00002b14
    x"00000000", -- 0x00002b18
    x"00000000", -- 0x00002b1c
    x"00000000", -- 0x00002b20
    x"00000000", -- 0x00002b24
    x"00000000", -- 0x00002b28
    x"00000000", -- 0x00002b2c
    x"00000000", -- 0x00002b30
    x"00000000", -- 0x00002b34
    x"00000000", -- 0x00002b38
    x"00000000", -- 0x00002b3c
    x"00000000", -- 0x00002b40
    x"00000000", -- 0x00002b44
    x"00000000", -- 0x00002b48
    x"00000000", -- 0x00002b4c
    x"00000000", -- 0x00002b50
    x"00000000", -- 0x00002b54
    x"00000000", -- 0x00002b58
    x"00000000", -- 0x00002b5c
    x"00000000", -- 0x00002b60
    x"00000000", -- 0x00002b64
    x"00000000", -- 0x00002b68
    x"00000000", -- 0x00002b6c
    x"00000000", -- 0x00002b70
    x"00000000", -- 0x00002b74
    x"00000000", -- 0x00002b78
    x"00000000", -- 0x00002b7c
    x"00000000", -- 0x00002b80
    x"00000000", -- 0x00002b84
    x"00000000", -- 0x00002b88
    x"00000000", -- 0x00002b8c
    x"00000000", -- 0x00002b90
    x"00000000", -- 0x00002b94
    x"00000000", -- 0x00002b98
    x"00000000", -- 0x00002b9c
    x"00000000", -- 0x00002ba0
    x"00000000", -- 0x00002ba4
    x"00000000", -- 0x00002ba8
    x"00000000", -- 0x00002bac
    x"00000000", -- 0x00002bb0
    x"00000000", -- 0x00002bb4
    x"00000000", -- 0x00002bb8
    x"00000000", -- 0x00002bbc
    x"00000000", -- 0x00002bc0
    x"00000000", -- 0x00002bc4
    x"00000000", -- 0x00002bc8
    x"00000000", -- 0x00002bcc
    x"00000000", -- 0x00002bd0
    x"00000000", -- 0x00002bd4
    x"00000000", -- 0x00002bd8
    x"00000000", -- 0x00002bdc
    x"00000000", -- 0x00002be0
    x"00000000", -- 0x00002be4
    x"00000000", -- 0x00002be8
    x"00000000", -- 0x00002bec
    x"00000000", -- 0x00002bf0
    x"00000000", -- 0x00002bf4
    x"00000000", -- 0x00002bf8
    x"00000000", -- 0x00002bfc
    x"00000000", -- 0x00002c00
    x"00000000", -- 0x00002c04
    x"00000000", -- 0x00002c08
    x"00000000", -- 0x00002c0c
    x"00000000", -- 0x00002c10
    x"00000000", -- 0x00002c14
    x"00000000", -- 0x00002c18
    x"00000000", -- 0x00002c1c
    x"00000000", -- 0x00002c20
    x"00000000", -- 0x00002c24
    x"00000000", -- 0x00002c28
    x"00000000", -- 0x00002c2c
    x"00000000", -- 0x00002c30
    x"00000000", -- 0x00002c34
    x"00000000", -- 0x00002c38
    x"00000000", -- 0x00002c3c
    x"00000000", -- 0x00002c40
    x"00000000", -- 0x00002c44
    x"00000000", -- 0x00002c48
    x"00000000", -- 0x00002c4c
    x"00000000", -- 0x00002c50
    x"00000000", -- 0x00002c54
    x"00000000", -- 0x00002c58
    x"00000000", -- 0x00002c5c
    x"00000000", -- 0x00002c60
    x"00000000", -- 0x00002c64
    x"00000000", -- 0x00002c68
    x"00000000", -- 0x00002c6c
    x"00000000", -- 0x00002c70
    x"00000000", -- 0x00002c74
    x"00000000", -- 0x00002c78
    x"00000000", -- 0x00002c7c
    x"00000000", -- 0x00002c80
    x"00000000", -- 0x00002c84
    x"00000000", -- 0x00002c88
    x"00000000", -- 0x00002c8c
    x"00000000", -- 0x00002c90
    x"00000000", -- 0x00002c94
    x"00000000", -- 0x00002c98
    x"00000000", -- 0x00002c9c
    x"00000000", -- 0x00002ca0
    x"00000000", -- 0x00002ca4
    x"00000000", -- 0x00002ca8
    x"00000000", -- 0x00002cac
    x"00000000", -- 0x00002cb0
    x"00000000", -- 0x00002cb4
    x"00000000", -- 0x00002cb8
    x"00000000", -- 0x00002cbc
    x"00000000", -- 0x00002cc0
    x"00000000", -- 0x00002cc4
    x"00000000", -- 0x00002cc8
    x"00000000", -- 0x00002ccc
    x"00000000", -- 0x00002cd0
    x"00000000", -- 0x00002cd4
    x"00000000", -- 0x00002cd8
    x"00000000", -- 0x00002cdc
    x"00000000", -- 0x00002ce0
    x"00000000", -- 0x00002ce4
    x"00000000", -- 0x00002ce8
    x"00000000", -- 0x00002cec
    x"00000000", -- 0x00002cf0
    x"00000000", -- 0x00002cf4
    x"00000000", -- 0x00002cf8
    x"00000000", -- 0x00002cfc
    x"00000000", -- 0x00002d00
    x"00000000", -- 0x00002d04
    x"00000000", -- 0x00002d08
    x"00000000", -- 0x00002d0c
    x"00000000", -- 0x00002d10
    x"00000000", -- 0x00002d14
    x"00000000", -- 0x00002d18
    x"00000000", -- 0x00002d1c
    x"00000000", -- 0x00002d20
    x"00000000", -- 0x00002d24
    x"00000000", -- 0x00002d28
    x"00000000", -- 0x00002d2c
    x"00000000", -- 0x00002d30
    x"00000000", -- 0x00002d34
    x"00000000", -- 0x00002d38
    x"00000000", -- 0x00002d3c
    x"00000000", -- 0x00002d40
    x"00000000", -- 0x00002d44
    x"00000000", -- 0x00002d48
    x"00000000", -- 0x00002d4c
    x"00000000", -- 0x00002d50
    x"00000000", -- 0x00002d54
    x"00000000", -- 0x00002d58
    x"00000000", -- 0x00002d5c
    x"00000000", -- 0x00002d60
    x"00000000", -- 0x00002d64
    x"00000000", -- 0x00002d68
    x"00000000", -- 0x00002d6c
    x"00000000", -- 0x00002d70
    x"00000000", -- 0x00002d74
    x"00000000", -- 0x00002d78
    x"00000000", -- 0x00002d7c
    x"00000000", -- 0x00002d80
    x"00000000", -- 0x00002d84
    x"00000000", -- 0x00002d88
    x"00000000", -- 0x00002d8c
    x"00000000", -- 0x00002d90
    x"00000000", -- 0x00002d94
    x"00000000", -- 0x00002d98
    x"00000000", -- 0x00002d9c
    x"00000000", -- 0x00002da0
    x"00000000", -- 0x00002da4
    x"00000000", -- 0x00002da8
    x"00000000", -- 0x00002dac
    x"00000000", -- 0x00002db0
    x"00000000", -- 0x00002db4
    x"00000000", -- 0x00002db8
    x"00000000", -- 0x00002dbc
    x"00000000", -- 0x00002dc0
    x"00000000", -- 0x00002dc4
    x"00000000", -- 0x00002dc8
    x"00000000", -- 0x00002dcc
    x"00000000", -- 0x00002dd0
    x"00000000", -- 0x00002dd4
    x"00000000", -- 0x00002dd8
    x"00000000", -- 0x00002ddc
    x"00000000", -- 0x00002de0
    x"00000000", -- 0x00002de4
    x"00000000", -- 0x00002de8
    x"00000000", -- 0x00002dec
    x"00000000", -- 0x00002df0
    x"00000000", -- 0x00002df4
    x"00000000", -- 0x00002df8
    x"00000000", -- 0x00002dfc
    x"00000000", -- 0x00002e00
    x"00000000", -- 0x00002e04
    x"00000000", -- 0x00002e08
    x"00000000", -- 0x00002e0c
    x"00000000", -- 0x00002e10
    x"00000000", -- 0x00002e14
    x"00000000", -- 0x00002e18
    x"00000000", -- 0x00002e1c
    x"00000000", -- 0x00002e20
    x"00000000", -- 0x00002e24
    x"00000000", -- 0x00002e28
    x"00000000", -- 0x00002e2c
    x"00000000", -- 0x00002e30
    x"00000000", -- 0x00002e34
    x"00000000", -- 0x00002e38
    x"00000000", -- 0x00002e3c
    x"00000000", -- 0x00002e40
    x"00000000", -- 0x00002e44
    x"00000000", -- 0x00002e48
    x"00000000", -- 0x00002e4c
    x"00000000", -- 0x00002e50
    x"00000000", -- 0x00002e54
    x"00000000", -- 0x00002e58
    x"00000000", -- 0x00002e5c
    x"00000000", -- 0x00002e60
    x"00000000", -- 0x00002e64
    x"00000000", -- 0x00002e68
    x"00000000", -- 0x00002e6c
    x"00000000", -- 0x00002e70
    x"00000000", -- 0x00002e74
    x"00000000", -- 0x00002e78
    x"00000000", -- 0x00002e7c
    x"00000000", -- 0x00002e80
    x"00000000", -- 0x00002e84
    x"00000000", -- 0x00002e88
    x"00000000", -- 0x00002e8c
    x"00000000", -- 0x00002e90
    x"00000000", -- 0x00002e94
    x"00000000", -- 0x00002e98
    x"00000000", -- 0x00002e9c
    x"00000000", -- 0x00002ea0
    x"00000000", -- 0x00002ea4
    x"00000000", -- 0x00002ea8
    x"00000000", -- 0x00002eac
    x"00000000", -- 0x00002eb0
    x"00000000", -- 0x00002eb4
    x"00000000", -- 0x00002eb8
    x"00000000", -- 0x00002ebc
    x"00000000", -- 0x00002ec0
    x"00000000", -- 0x00002ec4
    x"00000000", -- 0x00002ec8
    x"00000000", -- 0x00002ecc
    x"00000000", -- 0x00002ed0
    x"00000000", -- 0x00002ed4
    x"00000000", -- 0x00002ed8
    x"00000000", -- 0x00002edc
    x"00000000", -- 0x00002ee0
    x"00000000", -- 0x00002ee4
    x"00000000", -- 0x00002ee8
    x"00000000", -- 0x00002eec
    x"00000000", -- 0x00002ef0
    x"00000000", -- 0x00002ef4
    x"00000000", -- 0x00002ef8
    x"00000000", -- 0x00002efc
    x"00000000", -- 0x00002f00
    x"00000000", -- 0x00002f04
    x"00000000", -- 0x00002f08
    x"00000000", -- 0x00002f0c
    x"00000000", -- 0x00002f10
    x"00000000", -- 0x00002f14
    x"00000000", -- 0x00002f18
    x"00000000", -- 0x00002f1c
    x"00000000", -- 0x00002f20
    x"00000000", -- 0x00002f24
    x"00000000", -- 0x00002f28
    x"00000000", -- 0x00002f2c
    x"00000000", -- 0x00002f30
    x"00000000", -- 0x00002f34
    x"00000000", -- 0x00002f38
    x"00000000", -- 0x00002f3c
    x"00000000", -- 0x00002f40
    x"00000000", -- 0x00002f44
    x"00000000", -- 0x00002f48
    x"00000000", -- 0x00002f4c
    x"00000000", -- 0x00002f50
    x"00000000", -- 0x00002f54
    x"00000000", -- 0x00002f58
    x"00000000", -- 0x00002f5c
    x"00000000", -- 0x00002f60
    x"00000000", -- 0x00002f64
    x"00000000", -- 0x00002f68
    x"00000000", -- 0x00002f6c
    x"00000000", -- 0x00002f70
    x"00000000", -- 0x00002f74
    x"00000000", -- 0x00002f78
    x"00000000", -- 0x00002f7c
    x"00000000", -- 0x00002f80
    x"00000000", -- 0x00002f84
    x"00000000", -- 0x00002f88
    x"00000000", -- 0x00002f8c
    x"00000000", -- 0x00002f90
    x"00000000", -- 0x00002f94
    x"00000000", -- 0x00002f98
    x"00000000", -- 0x00002f9c
    x"00000000", -- 0x00002fa0
    x"00000000", -- 0x00002fa4
    x"00000000", -- 0x00002fa8
    x"00000000", -- 0x00002fac
    x"00000000", -- 0x00002fb0
    x"00000000", -- 0x00002fb4
    x"00000000", -- 0x00002fb8
    x"00000000", -- 0x00002fbc
    x"00000000", -- 0x00002fc0
    x"00000000", -- 0x00002fc4
    x"00000000", -- 0x00002fc8
    x"00000000", -- 0x00002fcc
    x"00000000", -- 0x00002fd0
    x"00000000", -- 0x00002fd4
    x"00000000", -- 0x00002fd8
    x"00000000", -- 0x00002fdc
    x"00000000", -- 0x00002fe0
    x"00000000", -- 0x00002fe4
    x"00000000", -- 0x00002fe8
    x"00000000", -- 0x00002fec
    x"00000000", -- 0x00002ff0
    x"00000000", -- 0x00002ff4
    x"00000000", -- 0x00002ff8
    x"00000000", -- 0x00002ffc
    x"00000000", -- 0x00003000
    x"00000000", -- 0x00003004
    x"00000000", -- 0x00003008
    x"00000000", -- 0x0000300c
    x"00000000", -- 0x00003010
    x"00000000", -- 0x00003014
    x"00000000", -- 0x00003018
    x"00000000", -- 0x0000301c
    x"00000000", -- 0x00003020
    x"00000000", -- 0x00003024
    x"00000000", -- 0x00003028
    x"00000000", -- 0x0000302c
    x"00000000", -- 0x00003030
    x"00000000", -- 0x00003034
    x"00000000", -- 0x00003038
    x"00000000", -- 0x0000303c
    x"00000000", -- 0x00003040
    x"00000000", -- 0x00003044
    x"00000000", -- 0x00003048
    x"00000000", -- 0x0000304c
    x"00000000", -- 0x00003050
    x"00000000", -- 0x00003054
    x"00000000", -- 0x00003058
    x"00000000", -- 0x0000305c
    x"00000000", -- 0x00003060
    x"00000000", -- 0x00003064
    x"00000000", -- 0x00003068
    x"00000000", -- 0x0000306c
    x"00000000", -- 0x00003070
    x"00000000", -- 0x00003074
    x"00000000", -- 0x00003078
    x"00000000", -- 0x0000307c
    x"00000000", -- 0x00003080
    x"00000000", -- 0x00003084
    x"00000000", -- 0x00003088
    x"00000000", -- 0x0000308c
    x"00000000", -- 0x00003090
    x"00000000", -- 0x00003094
    x"00000000", -- 0x00003098
    x"00000000", -- 0x0000309c
    x"00000000", -- 0x000030a0
    x"00000000", -- 0x000030a4
    x"00000000", -- 0x000030a8
    x"00000000", -- 0x000030ac
    x"00000000", -- 0x000030b0
    x"00000000", -- 0x000030b4
    x"00000000", -- 0x000030b8
    x"00000000", -- 0x000030bc
    x"00000000", -- 0x000030c0
    x"00000000", -- 0x000030c4
    x"00000000", -- 0x000030c8
    x"00000000", -- 0x000030cc
    x"00000000", -- 0x000030d0
    x"00000000", -- 0x000030d4
    x"00000000", -- 0x000030d8
    x"00000000", -- 0x000030dc
    x"00000000", -- 0x000030e0
    x"00000000", -- 0x000030e4
    x"00000000", -- 0x000030e8
    x"00000000", -- 0x000030ec
    x"00000000", -- 0x000030f0
    x"00000000", -- 0x000030f4
    x"00000000", -- 0x000030f8
    x"00000000", -- 0x000030fc
    x"00000000", -- 0x00003100
    x"00000000", -- 0x00003104
    x"00000000", -- 0x00003108
    x"00000000", -- 0x0000310c
    x"00000000", -- 0x00003110
    x"00000000", -- 0x00003114
    x"00000000", -- 0x00003118
    x"00000000", -- 0x0000311c
    x"00000000", -- 0x00003120
    x"00000000", -- 0x00003124
    x"00000000", -- 0x00003128
    x"00000000", -- 0x0000312c
    x"00000000", -- 0x00003130
    x"00000000", -- 0x00003134
    x"00000000", -- 0x00003138
    x"00000000", -- 0x0000313c
    x"00000000", -- 0x00003140
    x"00000000", -- 0x00003144
    x"00000000", -- 0x00003148
    x"00000000", -- 0x0000314c
    x"00000000", -- 0x00003150
    x"00000000", -- 0x00003154
    x"00000000", -- 0x00003158
    x"00000000", -- 0x0000315c
    x"00000000", -- 0x00003160
    x"00000000", -- 0x00003164
    x"00000000", -- 0x00003168
    x"00000000", -- 0x0000316c
    x"00000000", -- 0x00003170
    x"00000000", -- 0x00003174
    x"00000000", -- 0x00003178
    x"00000000", -- 0x0000317c
    x"00000000", -- 0x00003180
    x"00000000", -- 0x00003184
    x"00000000", -- 0x00003188
    x"00000000", -- 0x0000318c
    x"00000000", -- 0x00003190
    x"00000000", -- 0x00003194
    x"00000000", -- 0x00003198
    x"00000000", -- 0x0000319c
    x"00000000", -- 0x000031a0
    x"00000000", -- 0x000031a4
    x"00000000", -- 0x000031a8
    x"00000000", -- 0x000031ac
    x"00000000", -- 0x000031b0
    x"00000000", -- 0x000031b4
    x"00000000", -- 0x000031b8
    x"00000000", -- 0x000031bc
    x"00000000", -- 0x000031c0
    x"00000000", -- 0x000031c4
    x"00000000", -- 0x000031c8
    x"00000000", -- 0x000031cc
    x"00000000", -- 0x000031d0
    x"00000000", -- 0x000031d4
    x"00000000", -- 0x000031d8
    x"00000000", -- 0x000031dc
    x"00000000", -- 0x000031e0
    x"00000000", -- 0x000031e4
    x"00000000", -- 0x000031e8
    x"00000000", -- 0x000031ec
    x"00000000", -- 0x000031f0
    x"00000000", -- 0x000031f4
    x"00000000", -- 0x000031f8
    x"00000000", -- 0x000031fc
    x"00000000", -- 0x00003200
    x"00000000", -- 0x00003204
    x"00000000", -- 0x00003208
    x"00000000", -- 0x0000320c
    x"00000000", -- 0x00003210
    x"00000000", -- 0x00003214
    x"00000000", -- 0x00003218
    x"00000000", -- 0x0000321c
    x"00000000", -- 0x00003220
    x"00000000", -- 0x00003224
    x"00000000", -- 0x00003228
    x"00000000", -- 0x0000322c
    x"00000000", -- 0x00003230
    x"00000000", -- 0x00003234
    x"00000000", -- 0x00003238
    x"00000000", -- 0x0000323c
    x"00000000", -- 0x00003240
    x"00000000", -- 0x00003244
    x"00000000", -- 0x00003248
    x"00000000", -- 0x0000324c
    x"00000000", -- 0x00003250
    x"00000000", -- 0x00003254
    x"00000000", -- 0x00003258
    x"00000000", -- 0x0000325c
    x"00000000", -- 0x00003260
    x"00000000", -- 0x00003264
    x"00000000", -- 0x00003268
    x"00000000", -- 0x0000326c
    x"00000000", -- 0x00003270
    x"00000000", -- 0x00003274
    x"00000000", -- 0x00003278
    x"00000000", -- 0x0000327c
    x"00000000", -- 0x00003280
    x"00000000", -- 0x00003284
    x"00000000", -- 0x00003288
    x"00000000", -- 0x0000328c
    x"00000000", -- 0x00003290
    x"00000000", -- 0x00003294
    x"00000000", -- 0x00003298
    x"00000000", -- 0x0000329c
    x"00000000", -- 0x000032a0
    x"00000000", -- 0x000032a4
    x"00000000", -- 0x000032a8
    x"00000000", -- 0x000032ac
    x"00000000", -- 0x000032b0
    x"00000000", -- 0x000032b4
    x"00000000", -- 0x000032b8
    x"00000000", -- 0x000032bc
    x"00000000", -- 0x000032c0
    x"00000000", -- 0x000032c4
    x"00000000", -- 0x000032c8
    x"00000000", -- 0x000032cc
    x"00000000", -- 0x000032d0
    x"00000000", -- 0x000032d4
    x"00000000", -- 0x000032d8
    x"00000000", -- 0x000032dc
    x"00000000", -- 0x000032e0
    x"00000000", -- 0x000032e4
    x"00000000", -- 0x000032e8
    x"00000000", -- 0x000032ec
    x"00000000", -- 0x000032f0
    x"00000000", -- 0x000032f4
    x"00000000", -- 0x000032f8
    x"00000000", -- 0x000032fc
    x"00000000", -- 0x00003300
    x"00000000", -- 0x00003304
    x"00000000", -- 0x00003308
    x"00000000", -- 0x0000330c
    x"00000000", -- 0x00003310
    x"00000000", -- 0x00003314
    x"00000000", -- 0x00003318
    x"00000000", -- 0x0000331c
    x"00000000", -- 0x00003320
    x"00000000", -- 0x00003324
    x"00000000", -- 0x00003328
    x"00000000", -- 0x0000332c
    x"00000000", -- 0x00003330
    x"00000000", -- 0x00003334
    x"00000000", -- 0x00003338
    x"00000000", -- 0x0000333c
    x"00000000", -- 0x00003340
    x"00000000", -- 0x00003344
    x"00000000", -- 0x00003348
    x"00000000", -- 0x0000334c
    x"00000000", -- 0x00003350
    x"00000000", -- 0x00003354
    x"00000000", -- 0x00003358
    x"00000000", -- 0x0000335c
    x"00000000", -- 0x00003360
    x"00000000", -- 0x00003364
    x"00000000", -- 0x00003368
    x"00000000", -- 0x0000336c
    x"00000000", -- 0x00003370
    x"00000000", -- 0x00003374
    x"00000000", -- 0x00003378
    x"00000000", -- 0x0000337c
    x"00000000", -- 0x00003380
    x"00000000", -- 0x00003384
    x"00000000", -- 0x00003388
    x"00000000", -- 0x0000338c
    x"00000000", -- 0x00003390
    x"00000000", -- 0x00003394
    x"00000000", -- 0x00003398
    x"00000000", -- 0x0000339c
    x"00000000", -- 0x000033a0
    x"00000000", -- 0x000033a4
    x"00000000", -- 0x000033a8
    x"00000000", -- 0x000033ac
    x"00000000", -- 0x000033b0
    x"00000000", -- 0x000033b4
    x"00000000", -- 0x000033b8
    x"00000000", -- 0x000033bc
    x"00000000", -- 0x000033c0
    x"00000000", -- 0x000033c4
    x"00000000", -- 0x000033c8
    x"00000000", -- 0x000033cc
    x"00000000", -- 0x000033d0
    x"00000000", -- 0x000033d4
    x"00000000", -- 0x000033d8
    x"00000000", -- 0x000033dc
    x"00000000", -- 0x000033e0
    x"00000000", -- 0x000033e4
    x"00000000", -- 0x000033e8
    x"00000000", -- 0x000033ec
    x"00000000", -- 0x000033f0
    x"00000000", -- 0x000033f4
    x"00000000", -- 0x000033f8
    x"00000000", -- 0x000033fc
    x"00000000", -- 0x00003400
    x"00000000", -- 0x00003404
    x"00000000", -- 0x00003408
    x"00000000", -- 0x0000340c
    x"00000000", -- 0x00003410
    x"00000000", -- 0x00003414
    x"00000000", -- 0x00003418
    x"00000000", -- 0x0000341c
    x"00000000", -- 0x00003420
    x"00000000", -- 0x00003424
    x"00000000", -- 0x00003428
    x"00000000", -- 0x0000342c
    x"00000000", -- 0x00003430
    x"00000000", -- 0x00003434
    x"00000000", -- 0x00003438
    x"00000000", -- 0x0000343c
    x"00000000", -- 0x00003440
    x"00000000", -- 0x00003444
    x"00000000", -- 0x00003448
    x"00000000", -- 0x0000344c
    x"00000000", -- 0x00003450
    x"00000000", -- 0x00003454
    x"00000000", -- 0x00003458
    x"00000000", -- 0x0000345c
    x"00000000", -- 0x00003460
    x"00000000", -- 0x00003464
    x"00000000", -- 0x00003468
    x"00000000", -- 0x0000346c
    x"00000000", -- 0x00003470
    x"00000000", -- 0x00003474
    x"00000000", -- 0x00003478
    x"00000000", -- 0x0000347c
    x"00000000", -- 0x00003480
    x"00000000", -- 0x00003484
    x"00000000", -- 0x00003488
    x"00000000", -- 0x0000348c
    x"00000000", -- 0x00003490
    x"00000000", -- 0x00003494
    x"00000000", -- 0x00003498
    x"00000000", -- 0x0000349c
    x"00000000", -- 0x000034a0
    x"00000000", -- 0x000034a4
    x"00000000", -- 0x000034a8
    x"00000000", -- 0x000034ac
    x"00000000", -- 0x000034b0
    x"00000000", -- 0x000034b4
    x"00000000", -- 0x000034b8
    x"00000000", -- 0x000034bc
    x"00000000", -- 0x000034c0
    x"00000000", -- 0x000034c4
    x"00000000", -- 0x000034c8
    x"00000000", -- 0x000034cc
    x"00000000", -- 0x000034d0
    x"00000000", -- 0x000034d4
    x"00000000", -- 0x000034d8
    x"00000000", -- 0x000034dc
    x"00000000", -- 0x000034e0
    x"00000000", -- 0x000034e4
    x"00000000", -- 0x000034e8
    x"00000000", -- 0x000034ec
    x"00000000", -- 0x000034f0
    x"00000000", -- 0x000034f4
    x"00000000", -- 0x000034f8
    x"00000000", -- 0x000034fc
    x"00000000", -- 0x00003500
    x"00000000", -- 0x00003504
    x"00000000", -- 0x00003508
    x"00000000", -- 0x0000350c
    x"00000000", -- 0x00003510
    x"00000000", -- 0x00003514
    x"00000000", -- 0x00003518
    x"00000000", -- 0x0000351c
    x"00000000", -- 0x00003520
    x"00000000", -- 0x00003524
    x"00000000", -- 0x00003528
    x"00000000", -- 0x0000352c
    x"00000000", -- 0x00003530
    x"00000000", -- 0x00003534
    x"00000000", -- 0x00003538
    x"00000000", -- 0x0000353c
    x"00000000", -- 0x00003540
    x"00000000", -- 0x00003544
    x"00000000", -- 0x00003548
    x"00000000", -- 0x0000354c
    x"00000000", -- 0x00003550
    x"00000000", -- 0x00003554
    x"00000000", -- 0x00003558
    x"00000000", -- 0x0000355c
    x"00000000", -- 0x00003560
    x"00000000", -- 0x00003564
    x"00000000", -- 0x00003568
    x"00000000", -- 0x0000356c
    x"00000000", -- 0x00003570
    x"00000000", -- 0x00003574
    x"00000000", -- 0x00003578
    x"00000000", -- 0x0000357c
    x"00000000", -- 0x00003580
    x"00000000", -- 0x00003584
    x"00000000", -- 0x00003588
    x"00000000", -- 0x0000358c
    x"00000000", -- 0x00003590
    x"00000000", -- 0x00003594
    x"00000000", -- 0x00003598
    x"00000000", -- 0x0000359c
    x"00000000", -- 0x000035a0
    x"00000000", -- 0x000035a4
    x"00000000", -- 0x000035a8
    x"00000000", -- 0x000035ac
    x"00000000", -- 0x000035b0
    x"00000000", -- 0x000035b4
    x"00000000", -- 0x000035b8
    x"00000000", -- 0x000035bc
    x"00000000", -- 0x000035c0
    x"00000000", -- 0x000035c4
    x"00000000", -- 0x000035c8
    x"00000000", -- 0x000035cc
    x"00000000", -- 0x000035d0
    x"00000000", -- 0x000035d4
    x"00000000", -- 0x000035d8
    x"00000000", -- 0x000035dc
    x"00000000", -- 0x000035e0
    x"00000000", -- 0x000035e4
    x"00000000", -- 0x000035e8
    x"00000000", -- 0x000035ec
    x"00000000", -- 0x000035f0
    x"00000000", -- 0x000035f4
    x"00000000", -- 0x000035f8
    x"00000000", -- 0x000035fc
    x"00000000", -- 0x00003600
    x"00000000", -- 0x00003604
    x"00000000", -- 0x00003608
    x"00000000", -- 0x0000360c
    x"00000000", -- 0x00003610
    x"00000000", -- 0x00003614
    x"00000000", -- 0x00003618
    x"00000000", -- 0x0000361c
    x"00000000", -- 0x00003620
    x"00000000", -- 0x00003624
    x"00000000", -- 0x00003628
    x"00000000", -- 0x0000362c
    x"00000000", -- 0x00003630
    x"00000000", -- 0x00003634
    x"00000000", -- 0x00003638
    x"00000000", -- 0x0000363c
    x"00000000", -- 0x00003640
    x"00000000", -- 0x00003644
    x"00000000", -- 0x00003648
    x"00000000", -- 0x0000364c
    x"00000000", -- 0x00003650
    x"00000000", -- 0x00003654
    x"00000000", -- 0x00003658
    x"00000000", -- 0x0000365c
    x"00000000", -- 0x00003660
    x"00000000", -- 0x00003664
    x"00000000", -- 0x00003668
    x"00000000", -- 0x0000366c
    x"00000000", -- 0x00003670
    x"00000000", -- 0x00003674
    x"00000000", -- 0x00003678
    x"00000000", -- 0x0000367c
    x"00000000", -- 0x00003680
    x"00000000", -- 0x00003684
    x"00000000", -- 0x00003688
    x"00000000", -- 0x0000368c
    x"00000000", -- 0x00003690
    x"00000000", -- 0x00003694
    x"00000000", -- 0x00003698
    x"00000000", -- 0x0000369c
    x"00000000", -- 0x000036a0
    x"00000000", -- 0x000036a4
    x"00000000", -- 0x000036a8
    x"00000000", -- 0x000036ac
    x"00000000", -- 0x000036b0
    x"00000000", -- 0x000036b4
    x"00000000", -- 0x000036b8
    x"00000000", -- 0x000036bc
    x"00000000", -- 0x000036c0
    x"00000000", -- 0x000036c4
    x"00000000", -- 0x000036c8
    x"00000000", -- 0x000036cc
    x"00000000", -- 0x000036d0
    x"00000000", -- 0x000036d4
    x"00000000", -- 0x000036d8
    x"00000000", -- 0x000036dc
    x"00000000", -- 0x000036e0
    x"00000000", -- 0x000036e4
    x"00000000", -- 0x000036e8
    x"00000000", -- 0x000036ec
    x"00000000", -- 0x000036f0
    x"00000000", -- 0x000036f4
    x"00000000", -- 0x000036f8
    x"00000000", -- 0x000036fc
    x"00000000", -- 0x00003700
    x"00000000", -- 0x00003704
    x"00000000", -- 0x00003708
    x"00000000", -- 0x0000370c
    x"00000000", -- 0x00003710
    x"00000000", -- 0x00003714
    x"00000000", -- 0x00003718
    x"00000000", -- 0x0000371c
    x"00000000", -- 0x00003720
    x"00000000", -- 0x00003724
    x"00000000", -- 0x00003728
    x"00000000", -- 0x0000372c
    x"00000000", -- 0x00003730
    x"00000000", -- 0x00003734
    x"00000000", -- 0x00003738
    x"00000000", -- 0x0000373c
    x"00000000", -- 0x00003740
    x"00000000", -- 0x00003744
    x"00000000", -- 0x00003748
    x"00000000", -- 0x0000374c
    x"00000000", -- 0x00003750
    x"00000000", -- 0x00003754
    x"00000000", -- 0x00003758
    x"00000000", -- 0x0000375c
    x"00000000", -- 0x00003760
    x"00000000", -- 0x00003764
    x"00000000", -- 0x00003768
    x"00000000", -- 0x0000376c
    x"00000000", -- 0x00003770
    x"00000000", -- 0x00003774
    x"00000000", -- 0x00003778
    x"00000000", -- 0x0000377c
    x"00000000", -- 0x00003780
    x"00000000", -- 0x00003784
    x"00000000", -- 0x00003788
    x"00000000", -- 0x0000378c
    x"00000000", -- 0x00003790
    x"00000000", -- 0x00003794
    x"00000000", -- 0x00003798
    x"00000000", -- 0x0000379c
    x"00000000", -- 0x000037a0
    x"00000000", -- 0x000037a4
    x"00000000", -- 0x000037a8
    x"00000000", -- 0x000037ac
    x"00000000", -- 0x000037b0
    x"00000000", -- 0x000037b4
    x"00000000", -- 0x000037b8
    x"00000000", -- 0x000037bc
    x"00000000", -- 0x000037c0
    x"00000000", -- 0x000037c4
    x"00000000", -- 0x000037c8
    x"00000000", -- 0x000037cc
    x"00000000", -- 0x000037d0
    x"00000000", -- 0x000037d4
    x"00000000", -- 0x000037d8
    x"00000000", -- 0x000037dc
    x"00000000", -- 0x000037e0
    x"00000000", -- 0x000037e4
    x"00000000", -- 0x000037e8
    x"00000000", -- 0x000037ec
    x"00000000", -- 0x000037f0
    x"00000000", -- 0x000037f4
    x"00000000", -- 0x000037f8
    x"00000000", -- 0x000037fc
    x"00000000", -- 0x00003800
    x"00000000", -- 0x00003804
    x"00000000", -- 0x00003808
    x"00000000", -- 0x0000380c
    x"00000000", -- 0x00003810
    x"00000000", -- 0x00003814
    x"00000000", -- 0x00003818
    x"00000000", -- 0x0000381c
    x"00000000", -- 0x00003820
    x"00000000", -- 0x00003824
    x"00000000", -- 0x00003828
    x"00000000", -- 0x0000382c
    x"00000000", -- 0x00003830
    x"00000000", -- 0x00003834
    x"00000000", -- 0x00003838
    x"00000000", -- 0x0000383c
    x"00000000", -- 0x00003840
    x"00000000", -- 0x00003844
    x"00000000", -- 0x00003848
    x"00000000", -- 0x0000384c
    x"00000000", -- 0x00003850
    x"00000000", -- 0x00003854
    x"00000000", -- 0x00003858
    x"00000000", -- 0x0000385c
    x"00000000", -- 0x00003860
    x"00000000", -- 0x00003864
    x"00000000", -- 0x00003868
    x"00000000", -- 0x0000386c
    x"00000000", -- 0x00003870
    x"00000000", -- 0x00003874
    x"00000000", -- 0x00003878
    x"00000000", -- 0x0000387c
    x"00000000", -- 0x00003880
    x"00000000", -- 0x00003884
    x"00000000", -- 0x00003888
    x"00000000", -- 0x0000388c
    x"00000000", -- 0x00003890
    x"00000000", -- 0x00003894
    x"00000000", -- 0x00003898
    x"00000000", -- 0x0000389c
    x"00000000", -- 0x000038a0
    x"00000000", -- 0x000038a4
    x"00000000", -- 0x000038a8
    x"00000000", -- 0x000038ac
    x"00000000", -- 0x000038b0
    x"00000000", -- 0x000038b4
    x"00000000", -- 0x000038b8
    x"00000000", -- 0x000038bc
    x"00000000", -- 0x000038c0
    x"00000000", -- 0x000038c4
    x"00000000", -- 0x000038c8
    x"00000000", -- 0x000038cc
    x"00000000", -- 0x000038d0
    x"00000000", -- 0x000038d4
    x"00000000", -- 0x000038d8
    x"00000000", -- 0x000038dc
    x"00000000", -- 0x000038e0
    x"00000000", -- 0x000038e4
    x"00000000", -- 0x000038e8
    x"00000000", -- 0x000038ec
    x"00000000", -- 0x000038f0
    x"00000000", -- 0x000038f4
    x"00000000", -- 0x000038f8
    x"00000000", -- 0x000038fc
    x"00000000", -- 0x00003900
    x"00000000", -- 0x00003904
    x"00000000", -- 0x00003908
    x"00000000", -- 0x0000390c
    x"00000000", -- 0x00003910
    x"00000000", -- 0x00003914
    x"00000000", -- 0x00003918
    x"00000000", -- 0x0000391c
    x"00000000", -- 0x00003920
    x"00000000", -- 0x00003924
    x"00000000", -- 0x00003928
    x"00000000", -- 0x0000392c
    x"00000000", -- 0x00003930
    x"00000000", -- 0x00003934
    x"00000000", -- 0x00003938
    x"00000000", -- 0x0000393c
    x"00000000", -- 0x00003940
    x"00000000", -- 0x00003944
    x"00000000", -- 0x00003948
    x"00000000", -- 0x0000394c
    x"00000000", -- 0x00003950
    x"00000000", -- 0x00003954
    x"00000000", -- 0x00003958
    x"00000000", -- 0x0000395c
    x"00000000", -- 0x00003960
    x"00000000", -- 0x00003964
    x"00000000", -- 0x00003968
    x"00000000", -- 0x0000396c
    x"00000000", -- 0x00003970
    x"00000000", -- 0x00003974
    x"00000000", -- 0x00003978
    x"00000000", -- 0x0000397c
    x"00000000", -- 0x00003980
    x"00000000", -- 0x00003984
    x"00000000", -- 0x00003988
    x"00000000", -- 0x0000398c
    x"00000000", -- 0x00003990
    x"00000000", -- 0x00003994
    x"00000000", -- 0x00003998
    x"00000000", -- 0x0000399c
    x"00000000", -- 0x000039a0
    x"00000000", -- 0x000039a4
    x"00000000", -- 0x000039a8
    x"00000000", -- 0x000039ac
    x"00000000", -- 0x000039b0
    x"00000000", -- 0x000039b4
    x"00000000", -- 0x000039b8
    x"00000000", -- 0x000039bc
    x"00000000", -- 0x000039c0
    x"00000000", -- 0x000039c4
    x"00000000", -- 0x000039c8
    x"00000000", -- 0x000039cc
    x"00000000", -- 0x000039d0
    x"00000000", -- 0x000039d4
    x"00000000", -- 0x000039d8
    x"00000000", -- 0x000039dc
    x"00000000", -- 0x000039e0
    x"00000000", -- 0x000039e4
    x"00000000", -- 0x000039e8
    x"00000000", -- 0x000039ec
    x"00000000", -- 0x000039f0
    x"00000000", -- 0x000039f4
    x"00000000", -- 0x000039f8
    x"00000000", -- 0x000039fc
    x"00000000", -- 0x00003a00
    x"00000000", -- 0x00003a04
    x"00000000", -- 0x00003a08
    x"00000000", -- 0x00003a0c
    x"00000000", -- 0x00003a10
    x"00000000", -- 0x00003a14
    x"00000000", -- 0x00003a18
    x"00000000", -- 0x00003a1c
    x"00000000", -- 0x00003a20
    x"00000000", -- 0x00003a24
    x"00000000", -- 0x00003a28
    x"00000000", -- 0x00003a2c
    x"00000000", -- 0x00003a30
    x"00000000", -- 0x00003a34
    x"00000000", -- 0x00003a38
    x"00000000", -- 0x00003a3c
    x"00000000", -- 0x00003a40
    x"00000000", -- 0x00003a44
    x"00000000", -- 0x00003a48
    x"00000000", -- 0x00003a4c
    x"00000000", -- 0x00003a50
    x"00000000", -- 0x00003a54
    x"00000000", -- 0x00003a58
    x"00000000", -- 0x00003a5c
    x"00000000", -- 0x00003a60
    x"00000000", -- 0x00003a64
    x"00000000", -- 0x00003a68
    x"00000000", -- 0x00003a6c
    x"00000000", -- 0x00003a70
    x"00000000", -- 0x00003a74
    x"00000000", -- 0x00003a78
    x"00000000", -- 0x00003a7c
    x"00000000", -- 0x00003a80
    x"00000000", -- 0x00003a84
    x"00000000", -- 0x00003a88
    x"00000000", -- 0x00003a8c
    x"00000000", -- 0x00003a90
    x"00000000", -- 0x00003a94
    x"00000000", -- 0x00003a98
    x"00000000", -- 0x00003a9c
    x"00000000", -- 0x00003aa0
    x"00000000", -- 0x00003aa4
    x"00000000", -- 0x00003aa8
    x"00000000", -- 0x00003aac
    x"00000000", -- 0x00003ab0
    x"00000000", -- 0x00003ab4
    x"00000000", -- 0x00003ab8
    x"00000000", -- 0x00003abc
    x"00000000", -- 0x00003ac0
    x"00000000", -- 0x00003ac4
    x"00000000", -- 0x00003ac8
    x"00000000", -- 0x00003acc
    x"00000000", -- 0x00003ad0
    x"00000000", -- 0x00003ad4
    x"00000000", -- 0x00003ad8
    x"00000000", -- 0x00003adc
    x"00000000", -- 0x00003ae0
    x"00000000", -- 0x00003ae4
    x"00000000", -- 0x00003ae8
    x"00000000", -- 0x00003aec
    x"00000000", -- 0x00003af0
    x"00000000", -- 0x00003af4
    x"00000000", -- 0x00003af8
    x"00000000", -- 0x00003afc
    x"00000000", -- 0x00003b00
    x"00000000", -- 0x00003b04
    x"00000000", -- 0x00003b08
    x"00000000", -- 0x00003b0c
    x"00000000", -- 0x00003b10
    x"00000000", -- 0x00003b14
    x"00000000", -- 0x00003b18
    x"00000000", -- 0x00003b1c
    x"00000000", -- 0x00003b20
    x"00000000", -- 0x00003b24
    x"00000000", -- 0x00003b28
    x"00000000", -- 0x00003b2c
    x"00000000", -- 0x00003b30
    x"00000000", -- 0x00003b34
    x"00000000", -- 0x00003b38
    x"00000000", -- 0x00003b3c
    x"00000000", -- 0x00003b40
    x"00000000", -- 0x00003b44
    x"00000000", -- 0x00003b48
    x"00000000", -- 0x00003b4c
    x"00000000", -- 0x00003b50
    x"00000000", -- 0x00003b54
    x"00000000", -- 0x00003b58
    x"00000000", -- 0x00003b5c
    x"00000000", -- 0x00003b60
    x"00000000", -- 0x00003b64
    x"00000000", -- 0x00003b68
    x"00000000", -- 0x00003b6c
    x"00000000", -- 0x00003b70
    x"00000000", -- 0x00003b74
    x"00000000", -- 0x00003b78
    x"00000000", -- 0x00003b7c
    x"00000000", -- 0x00003b80
    x"00000000", -- 0x00003b84
    x"00000000", -- 0x00003b88
    x"00000000", -- 0x00003b8c
    x"00000000", -- 0x00003b90
    x"00000000", -- 0x00003b94
    x"00000000", -- 0x00003b98
    x"00000000", -- 0x00003b9c
    x"00000000", -- 0x00003ba0
    x"00000000", -- 0x00003ba4
    x"00000000", -- 0x00003ba8
    x"00000000", -- 0x00003bac
    x"00000000", -- 0x00003bb0
    x"00000000", -- 0x00003bb4
    x"00000000", -- 0x00003bb8
    x"00000000", -- 0x00003bbc
    x"00000000", -- 0x00003bc0
    x"00000000", -- 0x00003bc4
    x"00000000", -- 0x00003bc8
    x"00000000", -- 0x00003bcc
    x"00000000", -- 0x00003bd0
    x"00000000", -- 0x00003bd4
    x"00000000", -- 0x00003bd8
    x"00000000", -- 0x00003bdc
    x"00000000", -- 0x00003be0
    x"00000000", -- 0x00003be4
    x"00000000", -- 0x00003be8
    x"00000000", -- 0x00003bec
    x"00000000", -- 0x00003bf0
    x"00000000", -- 0x00003bf4
    x"00000000", -- 0x00003bf8
    x"00000000", -- 0x00003bfc
    x"00000000", -- 0x00003c00
    x"00000000", -- 0x00003c04
    x"00000000", -- 0x00003c08
    x"00000000", -- 0x00003c0c
    x"00000000", -- 0x00003c10
    x"00000000", -- 0x00003c14
    x"00000000", -- 0x00003c18
    x"00000000", -- 0x00003c1c
    x"00000000", -- 0x00003c20
    x"00000000", -- 0x00003c24
    x"00000000", -- 0x00003c28
    x"00000000", -- 0x00003c2c
    x"00000000", -- 0x00003c30
    x"00000000", -- 0x00003c34
    x"00000000", -- 0x00003c38
    x"00000000", -- 0x00003c3c
    x"00000000", -- 0x00003c40
    x"00000000", -- 0x00003c44
    x"00000000", -- 0x00003c48
    x"00000000", -- 0x00003c4c
    x"00000000", -- 0x00003c50
    x"00000000", -- 0x00003c54
    x"00000000", -- 0x00003c58
    x"00000000", -- 0x00003c5c
    x"00000000", -- 0x00003c60
    x"00000000", -- 0x00003c64
    x"00000000", -- 0x00003c68
    x"00000000", -- 0x00003c6c
    x"00000000", -- 0x00003c70
    x"00000000", -- 0x00003c74
    x"00000000", -- 0x00003c78
    x"00000000", -- 0x00003c7c
    x"00000000", -- 0x00003c80
    x"00000000", -- 0x00003c84
    x"00000000", -- 0x00003c88
    x"00000000", -- 0x00003c8c
    x"00000000", -- 0x00003c90
    x"00000000", -- 0x00003c94
    x"00000000", -- 0x00003c98
    x"00000000", -- 0x00003c9c
    x"00000000", -- 0x00003ca0
    x"00000000", -- 0x00003ca4
    x"00000000", -- 0x00003ca8
    x"00000000", -- 0x00003cac
    x"00000000", -- 0x00003cb0
    x"00000000", -- 0x00003cb4
    x"00000000", -- 0x00003cb8
    x"00000000", -- 0x00003cbc
    x"00000000", -- 0x00003cc0
    x"00000000", -- 0x00003cc4
    x"00000000", -- 0x00003cc8
    x"00000000", -- 0x00003ccc
    x"00000000", -- 0x00003cd0
    x"00000000", -- 0x00003cd4
    x"00000000", -- 0x00003cd8
    x"00000000", -- 0x00003cdc
    x"00000000", -- 0x00003ce0
    x"00000000", -- 0x00003ce4
    x"00000000", -- 0x00003ce8
    x"00000000", -- 0x00003cec
    x"00000000", -- 0x00003cf0
    x"00000000", -- 0x00003cf4
    x"00000000", -- 0x00003cf8
    x"00000000", -- 0x00003cfc
    x"00000000", -- 0x00003d00
    x"00000000", -- 0x00003d04
    x"00000000", -- 0x00003d08
    x"00000000", -- 0x00003d0c
    x"00000000", -- 0x00003d10
    x"00000000", -- 0x00003d14
    x"00000000", -- 0x00003d18
    x"00000000", -- 0x00003d1c
    x"00000000", -- 0x00003d20
    x"00000000", -- 0x00003d24
    x"00000000", -- 0x00003d28
    x"00000000", -- 0x00003d2c
    x"00000000", -- 0x00003d30
    x"00000000", -- 0x00003d34
    x"00000000", -- 0x00003d38
    x"00000000", -- 0x00003d3c
    x"00000000", -- 0x00003d40
    x"00000000", -- 0x00003d44
    x"00000000", -- 0x00003d48
    x"00000000", -- 0x00003d4c
    x"00000000", -- 0x00003d50
    x"00000000", -- 0x00003d54
    x"00000000", -- 0x00003d58
    x"00000000", -- 0x00003d5c
    x"00000000", -- 0x00003d60
    x"00000000", -- 0x00003d64
    x"00000000", -- 0x00003d68
    x"00000000", -- 0x00003d6c
    x"00000000", -- 0x00003d70
    x"00000000", -- 0x00003d74
    x"00000000", -- 0x00003d78
    x"00000000", -- 0x00003d7c
    x"00000000", -- 0x00003d80
    x"00000000", -- 0x00003d84
    x"00000000", -- 0x00003d88
    x"00000000", -- 0x00003d8c
    x"00000000", -- 0x00003d90
    x"00000000", -- 0x00003d94
    x"00000000", -- 0x00003d98
    x"00000000", -- 0x00003d9c
    x"00000000", -- 0x00003da0
    x"00000000", -- 0x00003da4
    x"00000000", -- 0x00003da8
    x"00000000", -- 0x00003dac
    x"00000000", -- 0x00003db0
    x"00000000", -- 0x00003db4
    x"00000000", -- 0x00003db8
    x"00000000", -- 0x00003dbc
    x"00000000", -- 0x00003dc0
    x"00000000", -- 0x00003dc4
    x"00000000", -- 0x00003dc8
    x"00000000", -- 0x00003dcc
    x"00000000", -- 0x00003dd0
    x"00000000", -- 0x00003dd4
    x"00000000", -- 0x00003dd8
    x"00000000", -- 0x00003ddc
    x"00000000", -- 0x00003de0
    x"00000000", -- 0x00003de4
    x"00000000", -- 0x00003de8
    x"00000000", -- 0x00003dec
    x"00000000", -- 0x00003df0
    x"00000000", -- 0x00003df4
    x"00000000", -- 0x00003df8
    x"00000000", -- 0x00003dfc
    x"00000000", -- 0x00003e00
    x"00000000", -- 0x00003e04
    x"00000000", -- 0x00003e08
    x"00000000", -- 0x00003e0c
    x"00000000", -- 0x00003e10
    x"00000000", -- 0x00003e14
    x"00000000", -- 0x00003e18
    x"00000000", -- 0x00003e1c
    x"00000000", -- 0x00003e20
    x"00000000", -- 0x00003e24
    x"00000000", -- 0x00003e28
    x"00000000", -- 0x00003e2c
    x"00000000", -- 0x00003e30
    x"00000000", -- 0x00003e34
    x"00000000", -- 0x00003e38
    x"00000000", -- 0x00003e3c
    x"00000000", -- 0x00003e40
    x"00000000", -- 0x00003e44
    x"00000000", -- 0x00003e48
    x"00000000", -- 0x00003e4c
    x"00000000", -- 0x00003e50
    x"00000000", -- 0x00003e54
    x"00000000", -- 0x00003e58
    x"00000000", -- 0x00003e5c
    x"00000000", -- 0x00003e60
    x"00000000", -- 0x00003e64
    x"00000000", -- 0x00003e68
    x"00000000", -- 0x00003e6c
    x"00000000", -- 0x00003e70
    x"00000000", -- 0x00003e74
    x"00000000", -- 0x00003e78
    x"00000000", -- 0x00003e7c
    x"00000000", -- 0x00003e80
    x"00000000", -- 0x00003e84
    x"00000000", -- 0x00003e88
    x"00000000", -- 0x00003e8c
    x"00000000", -- 0x00003e90
    x"00000000", -- 0x00003e94
    x"00000000", -- 0x00003e98
    x"00000000", -- 0x00003e9c
    x"00000000", -- 0x00003ea0
    x"00000000", -- 0x00003ea4
    x"00000000", -- 0x00003ea8
    x"00000000", -- 0x00003eac
    x"00000000", -- 0x00003eb0
    x"00000000", -- 0x00003eb4
    x"00000000", -- 0x00003eb8
    x"00000000", -- 0x00003ebc
    x"00000000", -- 0x00003ec0
    x"00000000", -- 0x00003ec4
    x"00000000", -- 0x00003ec8
    x"00000000", -- 0x00003ecc
    x"00000000", -- 0x00003ed0
    x"00000000", -- 0x00003ed4
    x"00000000", -- 0x00003ed8
    x"00000000", -- 0x00003edc
    x"00000000", -- 0x00003ee0
    x"00000000", -- 0x00003ee4
    x"00000000", -- 0x00003ee8
    x"00000000", -- 0x00003eec
    x"00000000", -- 0x00003ef0
    x"00000000", -- 0x00003ef4
    x"00000000", -- 0x00003ef8
    x"00000000", -- 0x00003efc
    x"00000000", -- 0x00003f00
    x"00000000", -- 0x00003f04
    x"00000000", -- 0x00003f08
    x"00000000", -- 0x00003f0c
    x"00000000", -- 0x00003f10
    x"00000000", -- 0x00003f14
    x"00000000", -- 0x00003f18
    x"00000000", -- 0x00003f1c
    x"00000000", -- 0x00003f20
    x"00000000", -- 0x00003f24
    x"00000000", -- 0x00003f28
    x"00000000", -- 0x00003f2c
    x"00000000", -- 0x00003f30
    x"00000000", -- 0x00003f34
    x"00000000", -- 0x00003f38
    x"00000000", -- 0x00003f3c
    x"00000000", -- 0x00003f40
    x"00000000", -- 0x00003f44
    x"00000000", -- 0x00003f48
    x"00000000", -- 0x00003f4c
    x"00000000", -- 0x00003f50
    x"00000000", -- 0x00003f54
    x"00000000", -- 0x00003f58
    x"00000000", -- 0x00003f5c
    x"00000000", -- 0x00003f60
    x"00000000", -- 0x00003f64
    x"00000000", -- 0x00003f68
    x"00000000", -- 0x00003f6c
    x"00000000", -- 0x00003f70
    x"00000000", -- 0x00003f74
    x"00000000", -- 0x00003f78
    x"00000000", -- 0x00003f7c
    x"00000000", -- 0x00003f80
    x"00000000", -- 0x00003f84
    x"00000000", -- 0x00003f88
    x"00000000", -- 0x00003f8c
    x"00000000", -- 0x00003f90
    x"00000000", -- 0x00003f94
    x"00000000", -- 0x00003f98
    x"00000000", -- 0x00003f9c
    x"00000000", -- 0x00003fa0
    x"00000000", -- 0x00003fa4
    x"00000000", -- 0x00003fa8
    x"00000000", -- 0x00003fac
    x"00000000", -- 0x00003fb0
    x"00000000", -- 0x00003fb4
    x"00000000", -- 0x00003fb8
    x"00000000", -- 0x00003fbc
    x"00000000", -- 0x00003fc0
    x"00000000", -- 0x00003fc4
    x"00000000", -- 0x00003fc8
    x"00000000", -- 0x00003fcc
    x"00000000", -- 0x00003fd0
    x"00000000", -- 0x00003fd4
    x"00000000", -- 0x00003fd8
    x"00000000", -- 0x00003fdc
    x"00000000", -- 0x00003fe0
    x"00000000", -- 0x00003fe4
    x"00000000", -- 0x00003fe8
    x"00000000", -- 0x00003fec
    x"00000000", -- 0x00003ff0
    x"00000000", -- 0x00003ff4
    x"00000000", -- 0x00003ff8
    x"00000000"  -- 0x00003ffc
  );
begin
  ACK_O <= read_ack or write_ack;
  DAT_O <= DAT_O_i;

  write_ack <= STB_I and WE_I;

  lookup_proc: process(CLK_I)
    variable addr : integer range 0 to 2 ** (ADR_I'length - 2) - 1;
  begin
    if rising_edge(CLK_I) then
      read_ack <= '0';
      DAT_O_i  <= (others=>'-');

      if RST_I = '0' then            
        if STB_I = '1' then 

          if WE_I = '0' and read_ack = '0' then
            addr  := to_integer(unsigned(ADR_I(ADR_I'length - 1 downto 2)));
            DAT_O_i  <= memory(addr);
            read_ack <= '1';
          elsif WE_I = '1' then
            addr  := to_integer(unsigned(ADR_I(ADR_I'length - 1 downto 2)));
            for i in 3 downto 0 loop
              if SEL_I(i) = '1' then
                memory(addr)(8 * i + 7 downto 8 * i) <= DAT_I(8 * i + 7 downto 8 * i);
              end if;
            end loop;
          end if;
        end if;
      end if;
    end if;
  end process;
end architecture;