library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity {entity} is
 port(
  CLK_I  : in  std_logic;
  RST_I  : in  std_logic;
  STB_I  : in  std_logic;
  WE_I   : in  std_logic;
  SEL_I  : in  std_logic_vector(3 downto 0);
  ADR_I  : in  std_logic_vector(13 downto 0);
  DAT_I  : in  std_logic_vector(31 downto 0);
  DAT_O  : out std_logic_vector(31 downto 0);
  ACK_O  : out std_logic
  );
end entity;

architecture behavioral of {entity} is
  type memory_t is array (0 to 2 ** (ADR_I'length - 2) - 1) of std_logic_vector(31 downto 0);

  signal read_ack  : std_logic := '0';
  signal write_ack : std_logic;
  signal DAT_O_i   : std_logic_vector(31 downto 0) := (others=>'-');
  signal memory    : memory_t := (
    x"{code[0x00000003-0x00000000,1]}", -- 0x00000000
    x"{code[0x00000007-0x00000004,1]}", -- 0x00000004
    x"{code[0x0000000b-0x00000008,1]}", -- 0x00000008
    x"{code[0x0000000f-0x0000000c,1]}", -- 0x0000000c
    x"{code[0x00000013-0x00000010,1]}", -- 0x00000010
    x"{code[0x00000017-0x00000014,1]}", -- 0x00000014
    x"{code[0x0000001b-0x00000018,1]}", -- 0x00000018
    x"{code[0x0000001f-0x0000001c,1]}", -- 0x0000001c
    x"{code[0x00000023-0x00000020,1]}", -- 0x00000020
    x"{code[0x00000027-0x00000024,1]}", -- 0x00000024
    x"{code[0x0000002b-0x00000028,1]}", -- 0x00000028
    x"{code[0x0000002f-0x0000002c,1]}", -- 0x0000002c
    x"{code[0x00000033-0x00000030,1]}", -- 0x00000030
    x"{code[0x00000037-0x00000034,1]}", -- 0x00000034
    x"{code[0x0000003b-0x00000038,1]}", -- 0x00000038
    x"{code[0x0000003f-0x0000003c,1]}", -- 0x0000003c
    x"{code[0x00000043-0x00000040,1]}", -- 0x00000040
    x"{code[0x00000047-0x00000044,1]}", -- 0x00000044
    x"{code[0x0000004b-0x00000048,1]}", -- 0x00000048
    x"{code[0x0000004f-0x0000004c,1]}", -- 0x0000004c
    x"{code[0x00000053-0x00000050,1]}", -- 0x00000050
    x"{code[0x00000057-0x00000054,1]}", -- 0x00000054
    x"{code[0x0000005b-0x00000058,1]}", -- 0x00000058
    x"{code[0x0000005f-0x0000005c,1]}", -- 0x0000005c
    x"{code[0x00000063-0x00000060,1]}", -- 0x00000060
    x"{code[0x00000067-0x00000064,1]}", -- 0x00000064
    x"{code[0x0000006b-0x00000068,1]}", -- 0x00000068
    x"{code[0x0000006f-0x0000006c,1]}", -- 0x0000006c
    x"{code[0x00000073-0x00000070,1]}", -- 0x00000070
    x"{code[0x00000077-0x00000074,1]}", -- 0x00000074
    x"{code[0x0000007b-0x00000078,1]}", -- 0x00000078
    x"{code[0x0000007f-0x0000007c,1]}", -- 0x0000007c
    x"{code[0x00000083-0x00000080,1]}", -- 0x00000080
    x"{code[0x00000087-0x00000084,1]}", -- 0x00000084
    x"{code[0x0000008b-0x00000088,1]}", -- 0x00000088
    x"{code[0x0000008f-0x0000008c,1]}", -- 0x0000008c
    x"{code[0x00000093-0x00000090,1]}", -- 0x00000090
    x"{code[0x00000097-0x00000094,1]}", -- 0x00000094
    x"{code[0x0000009b-0x00000098,1]}", -- 0x00000098
    x"{code[0x0000009f-0x0000009c,1]}", -- 0x0000009c
    x"{code[0x000000a3-0x000000a0,1]}", -- 0x000000a0
    x"{code[0x000000a7-0x000000a4,1]}", -- 0x000000a4
    x"{code[0x000000ab-0x000000a8,1]}", -- 0x000000a8
    x"{code[0x000000af-0x000000ac,1]}", -- 0x000000ac
    x"{code[0x000000b3-0x000000b0,1]}", -- 0x000000b0
    x"{code[0x000000b7-0x000000b4,1]}", -- 0x000000b4
    x"{code[0x000000bb-0x000000b8,1]}", -- 0x000000b8
    x"{code[0x000000bf-0x000000bc,1]}", -- 0x000000bc
    x"{code[0x000000c3-0x000000c0,1]}", -- 0x000000c0
    x"{code[0x000000c7-0x000000c4,1]}", -- 0x000000c4
    x"{code[0x000000cb-0x000000c8,1]}", -- 0x000000c8
    x"{code[0x000000cf-0x000000cc,1]}", -- 0x000000cc
    x"{code[0x000000d3-0x000000d0,1]}", -- 0x000000d0
    x"{code[0x000000d7-0x000000d4,1]}", -- 0x000000d4
    x"{code[0x000000db-0x000000d8,1]}", -- 0x000000d8
    x"{code[0x000000df-0x000000dc,1]}", -- 0x000000dc
    x"{code[0x000000e3-0x000000e0,1]}", -- 0x000000e0
    x"{code[0x000000e7-0x000000e4,1]}", -- 0x000000e4
    x"{code[0x000000eb-0x000000e8,1]}", -- 0x000000e8
    x"{code[0x000000ef-0x000000ec,1]}", -- 0x000000ec
    x"{code[0x000000f3-0x000000f0,1]}", -- 0x000000f0
    x"{code[0x000000f7-0x000000f4,1]}", -- 0x000000f4
    x"{code[0x000000fb-0x000000f8,1]}", -- 0x000000f8
    x"{code[0x000000ff-0x000000fc,1]}", -- 0x000000fc
    x"{code[0x00000103-0x00000100,1]}", -- 0x00000100
    x"{code[0x00000107-0x00000104,1]}", -- 0x00000104
    x"{code[0x0000010b-0x00000108,1]}", -- 0x00000108
    x"{code[0x0000010f-0x0000010c,1]}", -- 0x0000010c
    x"{code[0x00000113-0x00000110,1]}", -- 0x00000110
    x"{code[0x00000117-0x00000114,1]}", -- 0x00000114
    x"{code[0x0000011b-0x00000118,1]}", -- 0x00000118
    x"{code[0x0000011f-0x0000011c,1]}", -- 0x0000011c
    x"{code[0x00000123-0x00000120,1]}", -- 0x00000120
    x"{code[0x00000127-0x00000124,1]}", -- 0x00000124
    x"{code[0x0000012b-0x00000128,1]}", -- 0x00000128
    x"{code[0x0000012f-0x0000012c,1]}", -- 0x0000012c
    x"{code[0x00000133-0x00000130,1]}", -- 0x00000130
    x"{code[0x00000137-0x00000134,1]}", -- 0x00000134
    x"{code[0x0000013b-0x00000138,1]}", -- 0x00000138
    x"{code[0x0000013f-0x0000013c,1]}", -- 0x0000013c
    x"{code[0x00000143-0x00000140,1]}", -- 0x00000140
    x"{code[0x00000147-0x00000144,1]}", -- 0x00000144
    x"{code[0x0000014b-0x00000148,1]}", -- 0x00000148
    x"{code[0x0000014f-0x0000014c,1]}", -- 0x0000014c
    x"{code[0x00000153-0x00000150,1]}", -- 0x00000150
    x"{code[0x00000157-0x00000154,1]}", -- 0x00000154
    x"{code[0x0000015b-0x00000158,1]}", -- 0x00000158
    x"{code[0x0000015f-0x0000015c,1]}", -- 0x0000015c
    x"{code[0x00000163-0x00000160,1]}", -- 0x00000160
    x"{code[0x00000167-0x00000164,1]}", -- 0x00000164
    x"{code[0x0000016b-0x00000168,1]}", -- 0x00000168
    x"{code[0x0000016f-0x0000016c,1]}", -- 0x0000016c
    x"{code[0x00000173-0x00000170,1]}", -- 0x00000170
    x"{code[0x00000177-0x00000174,1]}", -- 0x00000174
    x"{code[0x0000017b-0x00000178,1]}", -- 0x00000178
    x"{code[0x0000017f-0x0000017c,1]}", -- 0x0000017c
    x"{code[0x00000183-0x00000180,1]}", -- 0x00000180
    x"{code[0x00000187-0x00000184,1]}", -- 0x00000184
    x"{code[0x0000018b-0x00000188,1]}", -- 0x00000188
    x"{code[0x0000018f-0x0000018c,1]}", -- 0x0000018c
    x"{code[0x00000193-0x00000190,1]}", -- 0x00000190
    x"{code[0x00000197-0x00000194,1]}", -- 0x00000194
    x"{code[0x0000019b-0x00000198,1]}", -- 0x00000198
    x"{code[0x0000019f-0x0000019c,1]}", -- 0x0000019c
    x"{code[0x000001a3-0x000001a0,1]}", -- 0x000001a0
    x"{code[0x000001a7-0x000001a4,1]}", -- 0x000001a4
    x"{code[0x000001ab-0x000001a8,1]}", -- 0x000001a8
    x"{code[0x000001af-0x000001ac,1]}", -- 0x000001ac
    x"{code[0x000001b3-0x000001b0,1]}", -- 0x000001b0
    x"{code[0x000001b7-0x000001b4,1]}", -- 0x000001b4
    x"{code[0x000001bb-0x000001b8,1]}", -- 0x000001b8
    x"{code[0x000001bf-0x000001bc,1]}", -- 0x000001bc
    x"{code[0x000001c3-0x000001c0,1]}", -- 0x000001c0
    x"{code[0x000001c7-0x000001c4,1]}", -- 0x000001c4
    x"{code[0x000001cb-0x000001c8,1]}", -- 0x000001c8
    x"{code[0x000001cf-0x000001cc,1]}", -- 0x000001cc
    x"{code[0x000001d3-0x000001d0,1]}", -- 0x000001d0
    x"{code[0x000001d7-0x000001d4,1]}", -- 0x000001d4
    x"{code[0x000001db-0x000001d8,1]}", -- 0x000001d8
    x"{code[0x000001df-0x000001dc,1]}", -- 0x000001dc
    x"{code[0x000001e3-0x000001e0,1]}", -- 0x000001e0
    x"{code[0x000001e7-0x000001e4,1]}", -- 0x000001e4
    x"{code[0x000001eb-0x000001e8,1]}", -- 0x000001e8
    x"{code[0x000001ef-0x000001ec,1]}", -- 0x000001ec
    x"{code[0x000001f3-0x000001f0,1]}", -- 0x000001f0
    x"{code[0x000001f7-0x000001f4,1]}", -- 0x000001f4
    x"{code[0x000001fb-0x000001f8,1]}", -- 0x000001f8
    x"{code[0x000001ff-0x000001fc,1]}", -- 0x000001fc
    x"{code[0x00000203-0x00000200,1]}", -- 0x00000200
    x"{code[0x00000207-0x00000204,1]}", -- 0x00000204
    x"{code[0x0000020b-0x00000208,1]}", -- 0x00000208
    x"{code[0x0000020f-0x0000020c,1]}", -- 0x0000020c
    x"{code[0x00000213-0x00000210,1]}", -- 0x00000210
    x"{code[0x00000217-0x00000214,1]}", -- 0x00000214
    x"{code[0x0000021b-0x00000218,1]}", -- 0x00000218
    x"{code[0x0000021f-0x0000021c,1]}", -- 0x0000021c
    x"{code[0x00000223-0x00000220,1]}", -- 0x00000220
    x"{code[0x00000227-0x00000224,1]}", -- 0x00000224
    x"{code[0x0000022b-0x00000228,1]}", -- 0x00000228
    x"{code[0x0000022f-0x0000022c,1]}", -- 0x0000022c
    x"{code[0x00000233-0x00000230,1]}", -- 0x00000230
    x"{code[0x00000237-0x00000234,1]}", -- 0x00000234
    x"{code[0x0000023b-0x00000238,1]}", -- 0x00000238
    x"{code[0x0000023f-0x0000023c,1]}", -- 0x0000023c
    x"{code[0x00000243-0x00000240,1]}", -- 0x00000240
    x"{code[0x00000247-0x00000244,1]}", -- 0x00000244
    x"{code[0x0000024b-0x00000248,1]}", -- 0x00000248
    x"{code[0x0000024f-0x0000024c,1]}", -- 0x0000024c
    x"{code[0x00000253-0x00000250,1]}", -- 0x00000250
    x"{code[0x00000257-0x00000254,1]}", -- 0x00000254
    x"{code[0x0000025b-0x00000258,1]}", -- 0x00000258
    x"{code[0x0000025f-0x0000025c,1]}", -- 0x0000025c
    x"{code[0x00000263-0x00000260,1]}", -- 0x00000260
    x"{code[0x00000267-0x00000264,1]}", -- 0x00000264
    x"{code[0x0000026b-0x00000268,1]}", -- 0x00000268
    x"{code[0x0000026f-0x0000026c,1]}", -- 0x0000026c
    x"{code[0x00000273-0x00000270,1]}", -- 0x00000270
    x"{code[0x00000277-0x00000274,1]}", -- 0x00000274
    x"{code[0x0000027b-0x00000278,1]}", -- 0x00000278
    x"{code[0x0000027f-0x0000027c,1]}", -- 0x0000027c
    x"{code[0x00000283-0x00000280,1]}", -- 0x00000280
    x"{code[0x00000287-0x00000284,1]}", -- 0x00000284
    x"{code[0x0000028b-0x00000288,1]}", -- 0x00000288
    x"{code[0x0000028f-0x0000028c,1]}", -- 0x0000028c
    x"{code[0x00000293-0x00000290,1]}", -- 0x00000290
    x"{code[0x00000297-0x00000294,1]}", -- 0x00000294
    x"{code[0x0000029b-0x00000298,1]}", -- 0x00000298
    x"{code[0x0000029f-0x0000029c,1]}", -- 0x0000029c
    x"{code[0x000002a3-0x000002a0,1]}", -- 0x000002a0
    x"{code[0x000002a7-0x000002a4,1]}", -- 0x000002a4
    x"{code[0x000002ab-0x000002a8,1]}", -- 0x000002a8
    x"{code[0x000002af-0x000002ac,1]}", -- 0x000002ac
    x"{code[0x000002b3-0x000002b0,1]}", -- 0x000002b0
    x"{code[0x000002b7-0x000002b4,1]}", -- 0x000002b4
    x"{code[0x000002bb-0x000002b8,1]}", -- 0x000002b8
    x"{code[0x000002bf-0x000002bc,1]}", -- 0x000002bc
    x"{code[0x000002c3-0x000002c0,1]}", -- 0x000002c0
    x"{code[0x000002c7-0x000002c4,1]}", -- 0x000002c4
    x"{code[0x000002cb-0x000002c8,1]}", -- 0x000002c8
    x"{code[0x000002cf-0x000002cc,1]}", -- 0x000002cc
    x"{code[0x000002d3-0x000002d0,1]}", -- 0x000002d0
    x"{code[0x000002d7-0x000002d4,1]}", -- 0x000002d4
    x"{code[0x000002db-0x000002d8,1]}", -- 0x000002d8
    x"{code[0x000002df-0x000002dc,1]}", -- 0x000002dc
    x"{code[0x000002e3-0x000002e0,1]}", -- 0x000002e0
    x"{code[0x000002e7-0x000002e4,1]}", -- 0x000002e4
    x"{code[0x000002eb-0x000002e8,1]}", -- 0x000002e8
    x"{code[0x000002ef-0x000002ec,1]}", -- 0x000002ec
    x"{code[0x000002f3-0x000002f0,1]}", -- 0x000002f0
    x"{code[0x000002f7-0x000002f4,1]}", -- 0x000002f4
    x"{code[0x000002fb-0x000002f8,1]}", -- 0x000002f8
    x"{code[0x000002ff-0x000002fc,1]}", -- 0x000002fc
    x"{code[0x00000303-0x00000300,1]}", -- 0x00000300
    x"{code[0x00000307-0x00000304,1]}", -- 0x00000304
    x"{code[0x0000030b-0x00000308,1]}", -- 0x00000308
    x"{code[0x0000030f-0x0000030c,1]}", -- 0x0000030c
    x"{code[0x00000313-0x00000310,1]}", -- 0x00000310
    x"{code[0x00000317-0x00000314,1]}", -- 0x00000314
    x"{code[0x0000031b-0x00000318,1]}", -- 0x00000318
    x"{code[0x0000031f-0x0000031c,1]}", -- 0x0000031c
    x"{code[0x00000323-0x00000320,1]}", -- 0x00000320
    x"{code[0x00000327-0x00000324,1]}", -- 0x00000324
    x"{code[0x0000032b-0x00000328,1]}", -- 0x00000328
    x"{code[0x0000032f-0x0000032c,1]}", -- 0x0000032c
    x"{code[0x00000333-0x00000330,1]}", -- 0x00000330
    x"{code[0x00000337-0x00000334,1]}", -- 0x00000334
    x"{code[0x0000033b-0x00000338,1]}", -- 0x00000338
    x"{code[0x0000033f-0x0000033c,1]}", -- 0x0000033c
    x"{code[0x00000343-0x00000340,1]}", -- 0x00000340
    x"{code[0x00000347-0x00000344,1]}", -- 0x00000344
    x"{code[0x0000034b-0x00000348,1]}", -- 0x00000348
    x"{code[0x0000034f-0x0000034c,1]}", -- 0x0000034c
    x"{code[0x00000353-0x00000350,1]}", -- 0x00000350
    x"{code[0x00000357-0x00000354,1]}", -- 0x00000354
    x"{code[0x0000035b-0x00000358,1]}", -- 0x00000358
    x"{code[0x0000035f-0x0000035c,1]}", -- 0x0000035c
    x"{code[0x00000363-0x00000360,1]}", -- 0x00000360
    x"{code[0x00000367-0x00000364,1]}", -- 0x00000364
    x"{code[0x0000036b-0x00000368,1]}", -- 0x00000368
    x"{code[0x0000036f-0x0000036c,1]}", -- 0x0000036c
    x"{code[0x00000373-0x00000370,1]}", -- 0x00000370
    x"{code[0x00000377-0x00000374,1]}", -- 0x00000374
    x"{code[0x0000037b-0x00000378,1]}", -- 0x00000378
    x"{code[0x0000037f-0x0000037c,1]}", -- 0x0000037c
    x"{code[0x00000383-0x00000380,1]}", -- 0x00000380
    x"{code[0x00000387-0x00000384,1]}", -- 0x00000384
    x"{code[0x0000038b-0x00000388,1]}", -- 0x00000388
    x"{code[0x0000038f-0x0000038c,1]}", -- 0x0000038c
    x"{code[0x00000393-0x00000390,1]}", -- 0x00000390
    x"{code[0x00000397-0x00000394,1]}", -- 0x00000394
    x"{code[0x0000039b-0x00000398,1]}", -- 0x00000398
    x"{code[0x0000039f-0x0000039c,1]}", -- 0x0000039c
    x"{code[0x000003a3-0x000003a0,1]}", -- 0x000003a0
    x"{code[0x000003a7-0x000003a4,1]}", -- 0x000003a4
    x"{code[0x000003ab-0x000003a8,1]}", -- 0x000003a8
    x"{code[0x000003af-0x000003ac,1]}", -- 0x000003ac
    x"{code[0x000003b3-0x000003b0,1]}", -- 0x000003b0
    x"{code[0x000003b7-0x000003b4,1]}", -- 0x000003b4
    x"{code[0x000003bb-0x000003b8,1]}", -- 0x000003b8
    x"{code[0x000003bf-0x000003bc,1]}", -- 0x000003bc
    x"{code[0x000003c3-0x000003c0,1]}", -- 0x000003c0
    x"{code[0x000003c7-0x000003c4,1]}", -- 0x000003c4
    x"{code[0x000003cb-0x000003c8,1]}", -- 0x000003c8
    x"{code[0x000003cf-0x000003cc,1]}", -- 0x000003cc
    x"{code[0x000003d3-0x000003d0,1]}", -- 0x000003d0
    x"{code[0x000003d7-0x000003d4,1]}", -- 0x000003d4
    x"{code[0x000003db-0x000003d8,1]}", -- 0x000003d8
    x"{code[0x000003df-0x000003dc,1]}", -- 0x000003dc
    x"{code[0x000003e3-0x000003e0,1]}", -- 0x000003e0
    x"{code[0x000003e7-0x000003e4,1]}", -- 0x000003e4
    x"{code[0x000003eb-0x000003e8,1]}", -- 0x000003e8
    x"{code[0x000003ef-0x000003ec,1]}", -- 0x000003ec
    x"{code[0x000003f3-0x000003f0,1]}", -- 0x000003f0
    x"{code[0x000003f7-0x000003f4,1]}", -- 0x000003f4
    x"{code[0x000003fb-0x000003f8,1]}", -- 0x000003f8
    x"{code[0x000003ff-0x000003fc,1]}", -- 0x000003fc
    x"{code[0x00000403-0x00000400,1]}", -- 0x00000400
    x"{code[0x00000407-0x00000404,1]}", -- 0x00000404
    x"{code[0x0000040b-0x00000408,1]}", -- 0x00000408
    x"{code[0x0000040f-0x0000040c,1]}", -- 0x0000040c
    x"{code[0x00000413-0x00000410,1]}", -- 0x00000410
    x"{code[0x00000417-0x00000414,1]}", -- 0x00000414
    x"{code[0x0000041b-0x00000418,1]}", -- 0x00000418
    x"{code[0x0000041f-0x0000041c,1]}", -- 0x0000041c
    x"{code[0x00000423-0x00000420,1]}", -- 0x00000420
    x"{code[0x00000427-0x00000424,1]}", -- 0x00000424
    x"{code[0x0000042b-0x00000428,1]}", -- 0x00000428
    x"{code[0x0000042f-0x0000042c,1]}", -- 0x0000042c
    x"{code[0x00000433-0x00000430,1]}", -- 0x00000430
    x"{code[0x00000437-0x00000434,1]}", -- 0x00000434
    x"{code[0x0000043b-0x00000438,1]}", -- 0x00000438
    x"{code[0x0000043f-0x0000043c,1]}", -- 0x0000043c
    x"{code[0x00000443-0x00000440,1]}", -- 0x00000440
    x"{code[0x00000447-0x00000444,1]}", -- 0x00000444
    x"{code[0x0000044b-0x00000448,1]}", -- 0x00000448
    x"{code[0x0000044f-0x0000044c,1]}", -- 0x0000044c
    x"{code[0x00000453-0x00000450,1]}", -- 0x00000450
    x"{code[0x00000457-0x00000454,1]}", -- 0x00000454
    x"{code[0x0000045b-0x00000458,1]}", -- 0x00000458
    x"{code[0x0000045f-0x0000045c,1]}", -- 0x0000045c
    x"{code[0x00000463-0x00000460,1]}", -- 0x00000460
    x"{code[0x00000467-0x00000464,1]}", -- 0x00000464
    x"{code[0x0000046b-0x00000468,1]}", -- 0x00000468
    x"{code[0x0000046f-0x0000046c,1]}", -- 0x0000046c
    x"{code[0x00000473-0x00000470,1]}", -- 0x00000470
    x"{code[0x00000477-0x00000474,1]}", -- 0x00000474
    x"{code[0x0000047b-0x00000478,1]}", -- 0x00000478
    x"{code[0x0000047f-0x0000047c,1]}", -- 0x0000047c
    x"{code[0x00000483-0x00000480,1]}", -- 0x00000480
    x"{code[0x00000487-0x00000484,1]}", -- 0x00000484
    x"{code[0x0000048b-0x00000488,1]}", -- 0x00000488
    x"{code[0x0000048f-0x0000048c,1]}", -- 0x0000048c
    x"{code[0x00000493-0x00000490,1]}", -- 0x00000490
    x"{code[0x00000497-0x00000494,1]}", -- 0x00000494
    x"{code[0x0000049b-0x00000498,1]}", -- 0x00000498
    x"{code[0x0000049f-0x0000049c,1]}", -- 0x0000049c
    x"{code[0x000004a3-0x000004a0,1]}", -- 0x000004a0
    x"{code[0x000004a7-0x000004a4,1]}", -- 0x000004a4
    x"{code[0x000004ab-0x000004a8,1]}", -- 0x000004a8
    x"{code[0x000004af-0x000004ac,1]}", -- 0x000004ac
    x"{code[0x000004b3-0x000004b0,1]}", -- 0x000004b0
    x"{code[0x000004b7-0x000004b4,1]}", -- 0x000004b4
    x"{code[0x000004bb-0x000004b8,1]}", -- 0x000004b8
    x"{code[0x000004bf-0x000004bc,1]}", -- 0x000004bc
    x"{code[0x000004c3-0x000004c0,1]}", -- 0x000004c0
    x"{code[0x000004c7-0x000004c4,1]}", -- 0x000004c4
    x"{code[0x000004cb-0x000004c8,1]}", -- 0x000004c8
    x"{code[0x000004cf-0x000004cc,1]}", -- 0x000004cc
    x"{code[0x000004d3-0x000004d0,1]}", -- 0x000004d0
    x"{code[0x000004d7-0x000004d4,1]}", -- 0x000004d4
    x"{code[0x000004db-0x000004d8,1]}", -- 0x000004d8
    x"{code[0x000004df-0x000004dc,1]}", -- 0x000004dc
    x"{code[0x000004e3-0x000004e0,1]}", -- 0x000004e0
    x"{code[0x000004e7-0x000004e4,1]}", -- 0x000004e4
    x"{code[0x000004eb-0x000004e8,1]}", -- 0x000004e8
    x"{code[0x000004ef-0x000004ec,1]}", -- 0x000004ec
    x"{code[0x000004f3-0x000004f0,1]}", -- 0x000004f0
    x"{code[0x000004f7-0x000004f4,1]}", -- 0x000004f4
    x"{code[0x000004fb-0x000004f8,1]}", -- 0x000004f8
    x"{code[0x000004ff-0x000004fc,1]}", -- 0x000004fc
    x"{code[0x00000503-0x00000500,1]}", -- 0x00000500
    x"{code[0x00000507-0x00000504,1]}", -- 0x00000504
    x"{code[0x0000050b-0x00000508,1]}", -- 0x00000508
    x"{code[0x0000050f-0x0000050c,1]}", -- 0x0000050c
    x"{code[0x00000513-0x00000510,1]}", -- 0x00000510
    x"{code[0x00000517-0x00000514,1]}", -- 0x00000514
    x"{code[0x0000051b-0x00000518,1]}", -- 0x00000518
    x"{code[0x0000051f-0x0000051c,1]}", -- 0x0000051c
    x"{code[0x00000523-0x00000520,1]}", -- 0x00000520
    x"{code[0x00000527-0x00000524,1]}", -- 0x00000524
    x"{code[0x0000052b-0x00000528,1]}", -- 0x00000528
    x"{code[0x0000052f-0x0000052c,1]}", -- 0x0000052c
    x"{code[0x00000533-0x00000530,1]}", -- 0x00000530
    x"{code[0x00000537-0x00000534,1]}", -- 0x00000534
    x"{code[0x0000053b-0x00000538,1]}", -- 0x00000538
    x"{code[0x0000053f-0x0000053c,1]}", -- 0x0000053c
    x"{code[0x00000543-0x00000540,1]}", -- 0x00000540
    x"{code[0x00000547-0x00000544,1]}", -- 0x00000544
    x"{code[0x0000054b-0x00000548,1]}", -- 0x00000548
    x"{code[0x0000054f-0x0000054c,1]}", -- 0x0000054c
    x"{code[0x00000553-0x00000550,1]}", -- 0x00000550
    x"{code[0x00000557-0x00000554,1]}", -- 0x00000554
    x"{code[0x0000055b-0x00000558,1]}", -- 0x00000558
    x"{code[0x0000055f-0x0000055c,1]}", -- 0x0000055c
    x"{code[0x00000563-0x00000560,1]}", -- 0x00000560
    x"{code[0x00000567-0x00000564,1]}", -- 0x00000564
    x"{code[0x0000056b-0x00000568,1]}", -- 0x00000568
    x"{code[0x0000056f-0x0000056c,1]}", -- 0x0000056c
    x"{code[0x00000573-0x00000570,1]}", -- 0x00000570
    x"{code[0x00000577-0x00000574,1]}", -- 0x00000574
    x"{code[0x0000057b-0x00000578,1]}", -- 0x00000578
    x"{code[0x0000057f-0x0000057c,1]}", -- 0x0000057c
    x"{code[0x00000583-0x00000580,1]}", -- 0x00000580
    x"{code[0x00000587-0x00000584,1]}", -- 0x00000584
    x"{code[0x0000058b-0x00000588,1]}", -- 0x00000588
    x"{code[0x0000058f-0x0000058c,1]}", -- 0x0000058c
    x"{code[0x00000593-0x00000590,1]}", -- 0x00000590
    x"{code[0x00000597-0x00000594,1]}", -- 0x00000594
    x"{code[0x0000059b-0x00000598,1]}", -- 0x00000598
    x"{code[0x0000059f-0x0000059c,1]}", -- 0x0000059c
    x"{code[0x000005a3-0x000005a0,1]}", -- 0x000005a0
    x"{code[0x000005a7-0x000005a4,1]}", -- 0x000005a4
    x"{code[0x000005ab-0x000005a8,1]}", -- 0x000005a8
    x"{code[0x000005af-0x000005ac,1]}", -- 0x000005ac
    x"{code[0x000005b3-0x000005b0,1]}", -- 0x000005b0
    x"{code[0x000005b7-0x000005b4,1]}", -- 0x000005b4
    x"{code[0x000005bb-0x000005b8,1]}", -- 0x000005b8
    x"{code[0x000005bf-0x000005bc,1]}", -- 0x000005bc
    x"{code[0x000005c3-0x000005c0,1]}", -- 0x000005c0
    x"{code[0x000005c7-0x000005c4,1]}", -- 0x000005c4
    x"{code[0x000005cb-0x000005c8,1]}", -- 0x000005c8
    x"{code[0x000005cf-0x000005cc,1]}", -- 0x000005cc
    x"{code[0x000005d3-0x000005d0,1]}", -- 0x000005d0
    x"{code[0x000005d7-0x000005d4,1]}", -- 0x000005d4
    x"{code[0x000005db-0x000005d8,1]}", -- 0x000005d8
    x"{code[0x000005df-0x000005dc,1]}", -- 0x000005dc
    x"{code[0x000005e3-0x000005e0,1]}", -- 0x000005e0
    x"{code[0x000005e7-0x000005e4,1]}", -- 0x000005e4
    x"{code[0x000005eb-0x000005e8,1]}", -- 0x000005e8
    x"{code[0x000005ef-0x000005ec,1]}", -- 0x000005ec
    x"{code[0x000005f3-0x000005f0,1]}", -- 0x000005f0
    x"{code[0x000005f7-0x000005f4,1]}", -- 0x000005f4
    x"{code[0x000005fb-0x000005f8,1]}", -- 0x000005f8
    x"{code[0x000005ff-0x000005fc,1]}", -- 0x000005fc
    x"{code[0x00000603-0x00000600,1]}", -- 0x00000600
    x"{code[0x00000607-0x00000604,1]}", -- 0x00000604
    x"{code[0x0000060b-0x00000608,1]}", -- 0x00000608
    x"{code[0x0000060f-0x0000060c,1]}", -- 0x0000060c
    x"{code[0x00000613-0x00000610,1]}", -- 0x00000610
    x"{code[0x00000617-0x00000614,1]}", -- 0x00000614
    x"{code[0x0000061b-0x00000618,1]}", -- 0x00000618
    x"{code[0x0000061f-0x0000061c,1]}", -- 0x0000061c
    x"{code[0x00000623-0x00000620,1]}", -- 0x00000620
    x"{code[0x00000627-0x00000624,1]}", -- 0x00000624
    x"{code[0x0000062b-0x00000628,1]}", -- 0x00000628
    x"{code[0x0000062f-0x0000062c,1]}", -- 0x0000062c
    x"{code[0x00000633-0x00000630,1]}", -- 0x00000630
    x"{code[0x00000637-0x00000634,1]}", -- 0x00000634
    x"{code[0x0000063b-0x00000638,1]}", -- 0x00000638
    x"{code[0x0000063f-0x0000063c,1]}", -- 0x0000063c
    x"{code[0x00000643-0x00000640,1]}", -- 0x00000640
    x"{code[0x00000647-0x00000644,1]}", -- 0x00000644
    x"{code[0x0000064b-0x00000648,1]}", -- 0x00000648
    x"{code[0x0000064f-0x0000064c,1]}", -- 0x0000064c
    x"{code[0x00000653-0x00000650,1]}", -- 0x00000650
    x"{code[0x00000657-0x00000654,1]}", -- 0x00000654
    x"{code[0x0000065b-0x00000658,1]}", -- 0x00000658
    x"{code[0x0000065f-0x0000065c,1]}", -- 0x0000065c
    x"{code[0x00000663-0x00000660,1]}", -- 0x00000660
    x"{code[0x00000667-0x00000664,1]}", -- 0x00000664
    x"{code[0x0000066b-0x00000668,1]}", -- 0x00000668
    x"{code[0x0000066f-0x0000066c,1]}", -- 0x0000066c
    x"{code[0x00000673-0x00000670,1]}", -- 0x00000670
    x"{code[0x00000677-0x00000674,1]}", -- 0x00000674
    x"{code[0x0000067b-0x00000678,1]}", -- 0x00000678
    x"{code[0x0000067f-0x0000067c,1]}", -- 0x0000067c
    x"{code[0x00000683-0x00000680,1]}", -- 0x00000680
    x"{code[0x00000687-0x00000684,1]}", -- 0x00000684
    x"{code[0x0000068b-0x00000688,1]}", -- 0x00000688
    x"{code[0x0000068f-0x0000068c,1]}", -- 0x0000068c
    x"{code[0x00000693-0x00000690,1]}", -- 0x00000690
    x"{code[0x00000697-0x00000694,1]}", -- 0x00000694
    x"{code[0x0000069b-0x00000698,1]}", -- 0x00000698
    x"{code[0x0000069f-0x0000069c,1]}", -- 0x0000069c
    x"{code[0x000006a3-0x000006a0,1]}", -- 0x000006a0
    x"{code[0x000006a7-0x000006a4,1]}", -- 0x000006a4
    x"{code[0x000006ab-0x000006a8,1]}", -- 0x000006a8
    x"{code[0x000006af-0x000006ac,1]}", -- 0x000006ac
    x"{code[0x000006b3-0x000006b0,1]}", -- 0x000006b0
    x"{code[0x000006b7-0x000006b4,1]}", -- 0x000006b4
    x"{code[0x000006bb-0x000006b8,1]}", -- 0x000006b8
    x"{code[0x000006bf-0x000006bc,1]}", -- 0x000006bc
    x"{code[0x000006c3-0x000006c0,1]}", -- 0x000006c0
    x"{code[0x000006c7-0x000006c4,1]}", -- 0x000006c4
    x"{code[0x000006cb-0x000006c8,1]}", -- 0x000006c8
    x"{code[0x000006cf-0x000006cc,1]}", -- 0x000006cc
    x"{code[0x000006d3-0x000006d0,1]}", -- 0x000006d0
    x"{code[0x000006d7-0x000006d4,1]}", -- 0x000006d4
    x"{code[0x000006db-0x000006d8,1]}", -- 0x000006d8
    x"{code[0x000006df-0x000006dc,1]}", -- 0x000006dc
    x"{code[0x000006e3-0x000006e0,1]}", -- 0x000006e0
    x"{code[0x000006e7-0x000006e4,1]}", -- 0x000006e4
    x"{code[0x000006eb-0x000006e8,1]}", -- 0x000006e8
    x"{code[0x000006ef-0x000006ec,1]}", -- 0x000006ec
    x"{code[0x000006f3-0x000006f0,1]}", -- 0x000006f0
    x"{code[0x000006f7-0x000006f4,1]}", -- 0x000006f4
    x"{code[0x000006fb-0x000006f8,1]}", -- 0x000006f8
    x"{code[0x000006ff-0x000006fc,1]}", -- 0x000006fc
    x"{code[0x00000703-0x00000700,1]}", -- 0x00000700
    x"{code[0x00000707-0x00000704,1]}", -- 0x00000704
    x"{code[0x0000070b-0x00000708,1]}", -- 0x00000708
    x"{code[0x0000070f-0x0000070c,1]}", -- 0x0000070c
    x"{code[0x00000713-0x00000710,1]}", -- 0x00000710
    x"{code[0x00000717-0x00000714,1]}", -- 0x00000714
    x"{code[0x0000071b-0x00000718,1]}", -- 0x00000718
    x"{code[0x0000071f-0x0000071c,1]}", -- 0x0000071c
    x"{code[0x00000723-0x00000720,1]}", -- 0x00000720
    x"{code[0x00000727-0x00000724,1]}", -- 0x00000724
    x"{code[0x0000072b-0x00000728,1]}", -- 0x00000728
    x"{code[0x0000072f-0x0000072c,1]}", -- 0x0000072c
    x"{code[0x00000733-0x00000730,1]}", -- 0x00000730
    x"{code[0x00000737-0x00000734,1]}", -- 0x00000734
    x"{code[0x0000073b-0x00000738,1]}", -- 0x00000738
    x"{code[0x0000073f-0x0000073c,1]}", -- 0x0000073c
    x"{code[0x00000743-0x00000740,1]}", -- 0x00000740
    x"{code[0x00000747-0x00000744,1]}", -- 0x00000744
    x"{code[0x0000074b-0x00000748,1]}", -- 0x00000748
    x"{code[0x0000074f-0x0000074c,1]}", -- 0x0000074c
    x"{code[0x00000753-0x00000750,1]}", -- 0x00000750
    x"{code[0x00000757-0x00000754,1]}", -- 0x00000754
    x"{code[0x0000075b-0x00000758,1]}", -- 0x00000758
    x"{code[0x0000075f-0x0000075c,1]}", -- 0x0000075c
    x"{code[0x00000763-0x00000760,1]}", -- 0x00000760
    x"{code[0x00000767-0x00000764,1]}", -- 0x00000764
    x"{code[0x0000076b-0x00000768,1]}", -- 0x00000768
    x"{code[0x0000076f-0x0000076c,1]}", -- 0x0000076c
    x"{code[0x00000773-0x00000770,1]}", -- 0x00000770
    x"{code[0x00000777-0x00000774,1]}", -- 0x00000774
    x"{code[0x0000077b-0x00000778,1]}", -- 0x00000778
    x"{code[0x0000077f-0x0000077c,1]}", -- 0x0000077c
    x"{code[0x00000783-0x00000780,1]}", -- 0x00000780
    x"{code[0x00000787-0x00000784,1]}", -- 0x00000784
    x"{code[0x0000078b-0x00000788,1]}", -- 0x00000788
    x"{code[0x0000078f-0x0000078c,1]}", -- 0x0000078c
    x"{code[0x00000793-0x00000790,1]}", -- 0x00000790
    x"{code[0x00000797-0x00000794,1]}", -- 0x00000794
    x"{code[0x0000079b-0x00000798,1]}", -- 0x00000798
    x"{code[0x0000079f-0x0000079c,1]}", -- 0x0000079c
    x"{code[0x000007a3-0x000007a0,1]}", -- 0x000007a0
    x"{code[0x000007a7-0x000007a4,1]}", -- 0x000007a4
    x"{code[0x000007ab-0x000007a8,1]}", -- 0x000007a8
    x"{code[0x000007af-0x000007ac,1]}", -- 0x000007ac
    x"{code[0x000007b3-0x000007b0,1]}", -- 0x000007b0
    x"{code[0x000007b7-0x000007b4,1]}", -- 0x000007b4
    x"{code[0x000007bb-0x000007b8,1]}", -- 0x000007b8
    x"{code[0x000007bf-0x000007bc,1]}", -- 0x000007bc
    x"{code[0x000007c3-0x000007c0,1]}", -- 0x000007c0
    x"{code[0x000007c7-0x000007c4,1]}", -- 0x000007c4
    x"{code[0x000007cb-0x000007c8,1]}", -- 0x000007c8
    x"{code[0x000007cf-0x000007cc,1]}", -- 0x000007cc
    x"{code[0x000007d3-0x000007d0,1]}", -- 0x000007d0
    x"{code[0x000007d7-0x000007d4,1]}", -- 0x000007d4
    x"{code[0x000007db-0x000007d8,1]}", -- 0x000007d8
    x"{code[0x000007df-0x000007dc,1]}", -- 0x000007dc
    x"{code[0x000007e3-0x000007e0,1]}", -- 0x000007e0
    x"{code[0x000007e7-0x000007e4,1]}", -- 0x000007e4
    x"{code[0x000007eb-0x000007e8,1]}", -- 0x000007e8
    x"{code[0x000007ef-0x000007ec,1]}", -- 0x000007ec
    x"{code[0x000007f3-0x000007f0,1]}", -- 0x000007f0
    x"{code[0x000007f7-0x000007f4,1]}", -- 0x000007f4
    x"{code[0x000007fb-0x000007f8,1]}", -- 0x000007f8
    x"{code[0x000007ff-0x000007fc,1]}", -- 0x000007fc
    x"{code[0x00000803-0x00000800,1]}", -- 0x00000800
    x"{code[0x00000807-0x00000804,1]}", -- 0x00000804
    x"{code[0x0000080b-0x00000808,1]}", -- 0x00000808
    x"{code[0x0000080f-0x0000080c,1]}", -- 0x0000080c
    x"{code[0x00000813-0x00000810,1]}", -- 0x00000810
    x"{code[0x00000817-0x00000814,1]}", -- 0x00000814
    x"{code[0x0000081b-0x00000818,1]}", -- 0x00000818
    x"{code[0x0000081f-0x0000081c,1]}", -- 0x0000081c
    x"{code[0x00000823-0x00000820,1]}", -- 0x00000820
    x"{code[0x00000827-0x00000824,1]}", -- 0x00000824
    x"{code[0x0000082b-0x00000828,1]}", -- 0x00000828
    x"{code[0x0000082f-0x0000082c,1]}", -- 0x0000082c
    x"{code[0x00000833-0x00000830,1]}", -- 0x00000830
    x"{code[0x00000837-0x00000834,1]}", -- 0x00000834
    x"{code[0x0000083b-0x00000838,1]}", -- 0x00000838
    x"{code[0x0000083f-0x0000083c,1]}", -- 0x0000083c
    x"{code[0x00000843-0x00000840,1]}", -- 0x00000840
    x"{code[0x00000847-0x00000844,1]}", -- 0x00000844
    x"{code[0x0000084b-0x00000848,1]}", -- 0x00000848
    x"{code[0x0000084f-0x0000084c,1]}", -- 0x0000084c
    x"{code[0x00000853-0x00000850,1]}", -- 0x00000850
    x"{code[0x00000857-0x00000854,1]}", -- 0x00000854
    x"{code[0x0000085b-0x00000858,1]}", -- 0x00000858
    x"{code[0x0000085f-0x0000085c,1]}", -- 0x0000085c
    x"{code[0x00000863-0x00000860,1]}", -- 0x00000860
    x"{code[0x00000867-0x00000864,1]}", -- 0x00000864
    x"{code[0x0000086b-0x00000868,1]}", -- 0x00000868
    x"{code[0x0000086f-0x0000086c,1]}", -- 0x0000086c
    x"{code[0x00000873-0x00000870,1]}", -- 0x00000870
    x"{code[0x00000877-0x00000874,1]}", -- 0x00000874
    x"{code[0x0000087b-0x00000878,1]}", -- 0x00000878
    x"{code[0x0000087f-0x0000087c,1]}", -- 0x0000087c
    x"{code[0x00000883-0x00000880,1]}", -- 0x00000880
    x"{code[0x00000887-0x00000884,1]}", -- 0x00000884
    x"{code[0x0000088b-0x00000888,1]}", -- 0x00000888
    x"{code[0x0000088f-0x0000088c,1]}", -- 0x0000088c
    x"{code[0x00000893-0x00000890,1]}", -- 0x00000890
    x"{code[0x00000897-0x00000894,1]}", -- 0x00000894
    x"{code[0x0000089b-0x00000898,1]}", -- 0x00000898
    x"{code[0x0000089f-0x0000089c,1]}", -- 0x0000089c
    x"{code[0x000008a3-0x000008a0,1]}", -- 0x000008a0
    x"{code[0x000008a7-0x000008a4,1]}", -- 0x000008a4
    x"{code[0x000008ab-0x000008a8,1]}", -- 0x000008a8
    x"{code[0x000008af-0x000008ac,1]}", -- 0x000008ac
    x"{code[0x000008b3-0x000008b0,1]}", -- 0x000008b0
    x"{code[0x000008b7-0x000008b4,1]}", -- 0x000008b4
    x"{code[0x000008bb-0x000008b8,1]}", -- 0x000008b8
    x"{code[0x000008bf-0x000008bc,1]}", -- 0x000008bc
    x"{code[0x000008c3-0x000008c0,1]}", -- 0x000008c0
    x"{code[0x000008c7-0x000008c4,1]}", -- 0x000008c4
    x"{code[0x000008cb-0x000008c8,1]}", -- 0x000008c8
    x"{code[0x000008cf-0x000008cc,1]}", -- 0x000008cc
    x"{code[0x000008d3-0x000008d0,1]}", -- 0x000008d0
    x"{code[0x000008d7-0x000008d4,1]}", -- 0x000008d4
    x"{code[0x000008db-0x000008d8,1]}", -- 0x000008d8
    x"{code[0x000008df-0x000008dc,1]}", -- 0x000008dc
    x"{code[0x000008e3-0x000008e0,1]}", -- 0x000008e0
    x"{code[0x000008e7-0x000008e4,1]}", -- 0x000008e4
    x"{code[0x000008eb-0x000008e8,1]}", -- 0x000008e8
    x"{code[0x000008ef-0x000008ec,1]}", -- 0x000008ec
    x"{code[0x000008f3-0x000008f0,1]}", -- 0x000008f0
    x"{code[0x000008f7-0x000008f4,1]}", -- 0x000008f4
    x"{code[0x000008fb-0x000008f8,1]}", -- 0x000008f8
    x"{code[0x000008ff-0x000008fc,1]}", -- 0x000008fc
    x"{code[0x00000903-0x00000900,1]}", -- 0x00000900
    x"{code[0x00000907-0x00000904,1]}", -- 0x00000904
    x"{code[0x0000090b-0x00000908,1]}", -- 0x00000908
    x"{code[0x0000090f-0x0000090c,1]}", -- 0x0000090c
    x"{code[0x00000913-0x00000910,1]}", -- 0x00000910
    x"{code[0x00000917-0x00000914,1]}", -- 0x00000914
    x"{code[0x0000091b-0x00000918,1]}", -- 0x00000918
    x"{code[0x0000091f-0x0000091c,1]}", -- 0x0000091c
    x"{code[0x00000923-0x00000920,1]}", -- 0x00000920
    x"{code[0x00000927-0x00000924,1]}", -- 0x00000924
    x"{code[0x0000092b-0x00000928,1]}", -- 0x00000928
    x"{code[0x0000092f-0x0000092c,1]}", -- 0x0000092c
    x"{code[0x00000933-0x00000930,1]}", -- 0x00000930
    x"{code[0x00000937-0x00000934,1]}", -- 0x00000934
    x"{code[0x0000093b-0x00000938,1]}", -- 0x00000938
    x"{code[0x0000093f-0x0000093c,1]}", -- 0x0000093c
    x"{code[0x00000943-0x00000940,1]}", -- 0x00000940
    x"{code[0x00000947-0x00000944,1]}", -- 0x00000944
    x"{code[0x0000094b-0x00000948,1]}", -- 0x00000948
    x"{code[0x0000094f-0x0000094c,1]}", -- 0x0000094c
    x"{code[0x00000953-0x00000950,1]}", -- 0x00000950
    x"{code[0x00000957-0x00000954,1]}", -- 0x00000954
    x"{code[0x0000095b-0x00000958,1]}", -- 0x00000958
    x"{code[0x0000095f-0x0000095c,1]}", -- 0x0000095c
    x"{code[0x00000963-0x00000960,1]}", -- 0x00000960
    x"{code[0x00000967-0x00000964,1]}", -- 0x00000964
    x"{code[0x0000096b-0x00000968,1]}", -- 0x00000968
    x"{code[0x0000096f-0x0000096c,1]}", -- 0x0000096c
    x"{code[0x00000973-0x00000970,1]}", -- 0x00000970
    x"{code[0x00000977-0x00000974,1]}", -- 0x00000974
    x"{code[0x0000097b-0x00000978,1]}", -- 0x00000978
    x"{code[0x0000097f-0x0000097c,1]}", -- 0x0000097c
    x"{code[0x00000983-0x00000980,1]}", -- 0x00000980
    x"{code[0x00000987-0x00000984,1]}", -- 0x00000984
    x"{code[0x0000098b-0x00000988,1]}", -- 0x00000988
    x"{code[0x0000098f-0x0000098c,1]}", -- 0x0000098c
    x"{code[0x00000993-0x00000990,1]}", -- 0x00000990
    x"{code[0x00000997-0x00000994,1]}", -- 0x00000994
    x"{code[0x0000099b-0x00000998,1]}", -- 0x00000998
    x"{code[0x0000099f-0x0000099c,1]}", -- 0x0000099c
    x"{code[0x000009a3-0x000009a0,1]}", -- 0x000009a0
    x"{code[0x000009a7-0x000009a4,1]}", -- 0x000009a4
    x"{code[0x000009ab-0x000009a8,1]}", -- 0x000009a8
    x"{code[0x000009af-0x000009ac,1]}", -- 0x000009ac
    x"{code[0x000009b3-0x000009b0,1]}", -- 0x000009b0
    x"{code[0x000009b7-0x000009b4,1]}", -- 0x000009b4
    x"{code[0x000009bb-0x000009b8,1]}", -- 0x000009b8
    x"{code[0x000009bf-0x000009bc,1]}", -- 0x000009bc
    x"{code[0x000009c3-0x000009c0,1]}", -- 0x000009c0
    x"{code[0x000009c7-0x000009c4,1]}", -- 0x000009c4
    x"{code[0x000009cb-0x000009c8,1]}", -- 0x000009c8
    x"{code[0x000009cf-0x000009cc,1]}", -- 0x000009cc
    x"{code[0x000009d3-0x000009d0,1]}", -- 0x000009d0
    x"{code[0x000009d7-0x000009d4,1]}", -- 0x000009d4
    x"{code[0x000009db-0x000009d8,1]}", -- 0x000009d8
    x"{code[0x000009df-0x000009dc,1]}", -- 0x000009dc
    x"{code[0x000009e3-0x000009e0,1]}", -- 0x000009e0
    x"{code[0x000009e7-0x000009e4,1]}", -- 0x000009e4
    x"{code[0x000009eb-0x000009e8,1]}", -- 0x000009e8
    x"{code[0x000009ef-0x000009ec,1]}", -- 0x000009ec
    x"{code[0x000009f3-0x000009f0,1]}", -- 0x000009f0
    x"{code[0x000009f7-0x000009f4,1]}", -- 0x000009f4
    x"{code[0x000009fb-0x000009f8,1]}", -- 0x000009f8
    x"{code[0x000009ff-0x000009fc,1]}", -- 0x000009fc
    x"{code[0x00000a03-0x00000a00,1]}", -- 0x00000a00
    x"{code[0x00000a07-0x00000a04,1]}", -- 0x00000a04
    x"{code[0x00000a0b-0x00000a08,1]}", -- 0x00000a08
    x"{code[0x00000a0f-0x00000a0c,1]}", -- 0x00000a0c
    x"{code[0x00000a13-0x00000a10,1]}", -- 0x00000a10
    x"{code[0x00000a17-0x00000a14,1]}", -- 0x00000a14
    x"{code[0x00000a1b-0x00000a18,1]}", -- 0x00000a18
    x"{code[0x00000a1f-0x00000a1c,1]}", -- 0x00000a1c
    x"{code[0x00000a23-0x00000a20,1]}", -- 0x00000a20
    x"{code[0x00000a27-0x00000a24,1]}", -- 0x00000a24
    x"{code[0x00000a2b-0x00000a28,1]}", -- 0x00000a28
    x"{code[0x00000a2f-0x00000a2c,1]}", -- 0x00000a2c
    x"{code[0x00000a33-0x00000a30,1]}", -- 0x00000a30
    x"{code[0x00000a37-0x00000a34,1]}", -- 0x00000a34
    x"{code[0x00000a3b-0x00000a38,1]}", -- 0x00000a38
    x"{code[0x00000a3f-0x00000a3c,1]}", -- 0x00000a3c
    x"{code[0x00000a43-0x00000a40,1]}", -- 0x00000a40
    x"{code[0x00000a47-0x00000a44,1]}", -- 0x00000a44
    x"{code[0x00000a4b-0x00000a48,1]}", -- 0x00000a48
    x"{code[0x00000a4f-0x00000a4c,1]}", -- 0x00000a4c
    x"{code[0x00000a53-0x00000a50,1]}", -- 0x00000a50
    x"{code[0x00000a57-0x00000a54,1]}", -- 0x00000a54
    x"{code[0x00000a5b-0x00000a58,1]}", -- 0x00000a58
    x"{code[0x00000a5f-0x00000a5c,1]}", -- 0x00000a5c
    x"{code[0x00000a63-0x00000a60,1]}", -- 0x00000a60
    x"{code[0x00000a67-0x00000a64,1]}", -- 0x00000a64
    x"{code[0x00000a6b-0x00000a68,1]}", -- 0x00000a68
    x"{code[0x00000a6f-0x00000a6c,1]}", -- 0x00000a6c
    x"{code[0x00000a73-0x00000a70,1]}", -- 0x00000a70
    x"{code[0x00000a77-0x00000a74,1]}", -- 0x00000a74
    x"{code[0x00000a7b-0x00000a78,1]}", -- 0x00000a78
    x"{code[0x00000a7f-0x00000a7c,1]}", -- 0x00000a7c
    x"{code[0x00000a83-0x00000a80,1]}", -- 0x00000a80
    x"{code[0x00000a87-0x00000a84,1]}", -- 0x00000a84
    x"{code[0x00000a8b-0x00000a88,1]}", -- 0x00000a88
    x"{code[0x00000a8f-0x00000a8c,1]}", -- 0x00000a8c
    x"{code[0x00000a93-0x00000a90,1]}", -- 0x00000a90
    x"{code[0x00000a97-0x00000a94,1]}", -- 0x00000a94
    x"{code[0x00000a9b-0x00000a98,1]}", -- 0x00000a98
    x"{code[0x00000a9f-0x00000a9c,1]}", -- 0x00000a9c
    x"{code[0x00000aa3-0x00000aa0,1]}", -- 0x00000aa0
    x"{code[0x00000aa7-0x00000aa4,1]}", -- 0x00000aa4
    x"{code[0x00000aab-0x00000aa8,1]}", -- 0x00000aa8
    x"{code[0x00000aaf-0x00000aac,1]}", -- 0x00000aac
    x"{code[0x00000ab3-0x00000ab0,1]}", -- 0x00000ab0
    x"{code[0x00000ab7-0x00000ab4,1]}", -- 0x00000ab4
    x"{code[0x00000abb-0x00000ab8,1]}", -- 0x00000ab8
    x"{code[0x00000abf-0x00000abc,1]}", -- 0x00000abc
    x"{code[0x00000ac3-0x00000ac0,1]}", -- 0x00000ac0
    x"{code[0x00000ac7-0x00000ac4,1]}", -- 0x00000ac4
    x"{code[0x00000acb-0x00000ac8,1]}", -- 0x00000ac8
    x"{code[0x00000acf-0x00000acc,1]}", -- 0x00000acc
    x"{code[0x00000ad3-0x00000ad0,1]}", -- 0x00000ad0
    x"{code[0x00000ad7-0x00000ad4,1]}", -- 0x00000ad4
    x"{code[0x00000adb-0x00000ad8,1]}", -- 0x00000ad8
    x"{code[0x00000adf-0x00000adc,1]}", -- 0x00000adc
    x"{code[0x00000ae3-0x00000ae0,1]}", -- 0x00000ae0
    x"{code[0x00000ae7-0x00000ae4,1]}", -- 0x00000ae4
    x"{code[0x00000aeb-0x00000ae8,1]}", -- 0x00000ae8
    x"{code[0x00000aef-0x00000aec,1]}", -- 0x00000aec
    x"{code[0x00000af3-0x00000af0,1]}", -- 0x00000af0
    x"{code[0x00000af7-0x00000af4,1]}", -- 0x00000af4
    x"{code[0x00000afb-0x00000af8,1]}", -- 0x00000af8
    x"{code[0x00000aff-0x00000afc,1]}", -- 0x00000afc
    x"{code[0x00000b03-0x00000b00,1]}", -- 0x00000b00
    x"{code[0x00000b07-0x00000b04,1]}", -- 0x00000b04
    x"{code[0x00000b0b-0x00000b08,1]}", -- 0x00000b08
    x"{code[0x00000b0f-0x00000b0c,1]}", -- 0x00000b0c
    x"{code[0x00000b13-0x00000b10,1]}", -- 0x00000b10
    x"{code[0x00000b17-0x00000b14,1]}", -- 0x00000b14
    x"{code[0x00000b1b-0x00000b18,1]}", -- 0x00000b18
    x"{code[0x00000b1f-0x00000b1c,1]}", -- 0x00000b1c
    x"{code[0x00000b23-0x00000b20,1]}", -- 0x00000b20
    x"{code[0x00000b27-0x00000b24,1]}", -- 0x00000b24
    x"{code[0x00000b2b-0x00000b28,1]}", -- 0x00000b28
    x"{code[0x00000b2f-0x00000b2c,1]}", -- 0x00000b2c
    x"{code[0x00000b33-0x00000b30,1]}", -- 0x00000b30
    x"{code[0x00000b37-0x00000b34,1]}", -- 0x00000b34
    x"{code[0x00000b3b-0x00000b38,1]}", -- 0x00000b38
    x"{code[0x00000b3f-0x00000b3c,1]}", -- 0x00000b3c
    x"{code[0x00000b43-0x00000b40,1]}", -- 0x00000b40
    x"{code[0x00000b47-0x00000b44,1]}", -- 0x00000b44
    x"{code[0x00000b4b-0x00000b48,1]}", -- 0x00000b48
    x"{code[0x00000b4f-0x00000b4c,1]}", -- 0x00000b4c
    x"{code[0x00000b53-0x00000b50,1]}", -- 0x00000b50
    x"{code[0x00000b57-0x00000b54,1]}", -- 0x00000b54
    x"{code[0x00000b5b-0x00000b58,1]}", -- 0x00000b58
    x"{code[0x00000b5f-0x00000b5c,1]}", -- 0x00000b5c
    x"{code[0x00000b63-0x00000b60,1]}", -- 0x00000b60
    x"{code[0x00000b67-0x00000b64,1]}", -- 0x00000b64
    x"{code[0x00000b6b-0x00000b68,1]}", -- 0x00000b68
    x"{code[0x00000b6f-0x00000b6c,1]}", -- 0x00000b6c
    x"{code[0x00000b73-0x00000b70,1]}", -- 0x00000b70
    x"{code[0x00000b77-0x00000b74,1]}", -- 0x00000b74
    x"{code[0x00000b7b-0x00000b78,1]}", -- 0x00000b78
    x"{code[0x00000b7f-0x00000b7c,1]}", -- 0x00000b7c
    x"{code[0x00000b83-0x00000b80,1]}", -- 0x00000b80
    x"{code[0x00000b87-0x00000b84,1]}", -- 0x00000b84
    x"{code[0x00000b8b-0x00000b88,1]}", -- 0x00000b88
    x"{code[0x00000b8f-0x00000b8c,1]}", -- 0x00000b8c
    x"{code[0x00000b93-0x00000b90,1]}", -- 0x00000b90
    x"{code[0x00000b97-0x00000b94,1]}", -- 0x00000b94
    x"{code[0x00000b9b-0x00000b98,1]}", -- 0x00000b98
    x"{code[0x00000b9f-0x00000b9c,1]}", -- 0x00000b9c
    x"{code[0x00000ba3-0x00000ba0,1]}", -- 0x00000ba0
    x"{code[0x00000ba7-0x00000ba4,1]}", -- 0x00000ba4
    x"{code[0x00000bab-0x00000ba8,1]}", -- 0x00000ba8
    x"{code[0x00000baf-0x00000bac,1]}", -- 0x00000bac
    x"{code[0x00000bb3-0x00000bb0,1]}", -- 0x00000bb0
    x"{code[0x00000bb7-0x00000bb4,1]}", -- 0x00000bb4
    x"{code[0x00000bbb-0x00000bb8,1]}", -- 0x00000bb8
    x"{code[0x00000bbf-0x00000bbc,1]}", -- 0x00000bbc
    x"{code[0x00000bc3-0x00000bc0,1]}", -- 0x00000bc0
    x"{code[0x00000bc7-0x00000bc4,1]}", -- 0x00000bc4
    x"{code[0x00000bcb-0x00000bc8,1]}", -- 0x00000bc8
    x"{code[0x00000bcf-0x00000bcc,1]}", -- 0x00000bcc
    x"{code[0x00000bd3-0x00000bd0,1]}", -- 0x00000bd0
    x"{code[0x00000bd7-0x00000bd4,1]}", -- 0x00000bd4
    x"{code[0x00000bdb-0x00000bd8,1]}", -- 0x00000bd8
    x"{code[0x00000bdf-0x00000bdc,1]}", -- 0x00000bdc
    x"{code[0x00000be3-0x00000be0,1]}", -- 0x00000be0
    x"{code[0x00000be7-0x00000be4,1]}", -- 0x00000be4
    x"{code[0x00000beb-0x00000be8,1]}", -- 0x00000be8
    x"{code[0x00000bef-0x00000bec,1]}", -- 0x00000bec
    x"{code[0x00000bf3-0x00000bf0,1]}", -- 0x00000bf0
    x"{code[0x00000bf7-0x00000bf4,1]}", -- 0x00000bf4
    x"{code[0x00000bfb-0x00000bf8,1]}", -- 0x00000bf8
    x"{code[0x00000bff-0x00000bfc,1]}", -- 0x00000bfc
    x"{code[0x00000c03-0x00000c00,1]}", -- 0x00000c00
    x"{code[0x00000c07-0x00000c04,1]}", -- 0x00000c04
    x"{code[0x00000c0b-0x00000c08,1]}", -- 0x00000c08
    x"{code[0x00000c0f-0x00000c0c,1]}", -- 0x00000c0c
    x"{code[0x00000c13-0x00000c10,1]}", -- 0x00000c10
    x"{code[0x00000c17-0x00000c14,1]}", -- 0x00000c14
    x"{code[0x00000c1b-0x00000c18,1]}", -- 0x00000c18
    x"{code[0x00000c1f-0x00000c1c,1]}", -- 0x00000c1c
    x"{code[0x00000c23-0x00000c20,1]}", -- 0x00000c20
    x"{code[0x00000c27-0x00000c24,1]}", -- 0x00000c24
    x"{code[0x00000c2b-0x00000c28,1]}", -- 0x00000c28
    x"{code[0x00000c2f-0x00000c2c,1]}", -- 0x00000c2c
    x"{code[0x00000c33-0x00000c30,1]}", -- 0x00000c30
    x"{code[0x00000c37-0x00000c34,1]}", -- 0x00000c34
    x"{code[0x00000c3b-0x00000c38,1]}", -- 0x00000c38
    x"{code[0x00000c3f-0x00000c3c,1]}", -- 0x00000c3c
    x"{code[0x00000c43-0x00000c40,1]}", -- 0x00000c40
    x"{code[0x00000c47-0x00000c44,1]}", -- 0x00000c44
    x"{code[0x00000c4b-0x00000c48,1]}", -- 0x00000c48
    x"{code[0x00000c4f-0x00000c4c,1]}", -- 0x00000c4c
    x"{code[0x00000c53-0x00000c50,1]}", -- 0x00000c50
    x"{code[0x00000c57-0x00000c54,1]}", -- 0x00000c54
    x"{code[0x00000c5b-0x00000c58,1]}", -- 0x00000c58
    x"{code[0x00000c5f-0x00000c5c,1]}", -- 0x00000c5c
    x"{code[0x00000c63-0x00000c60,1]}", -- 0x00000c60
    x"{code[0x00000c67-0x00000c64,1]}", -- 0x00000c64
    x"{code[0x00000c6b-0x00000c68,1]}", -- 0x00000c68
    x"{code[0x00000c6f-0x00000c6c,1]}", -- 0x00000c6c
    x"{code[0x00000c73-0x00000c70,1]}", -- 0x00000c70
    x"{code[0x00000c77-0x00000c74,1]}", -- 0x00000c74
    x"{code[0x00000c7b-0x00000c78,1]}", -- 0x00000c78
    x"{code[0x00000c7f-0x00000c7c,1]}", -- 0x00000c7c
    x"{code[0x00000c83-0x00000c80,1]}", -- 0x00000c80
    x"{code[0x00000c87-0x00000c84,1]}", -- 0x00000c84
    x"{code[0x00000c8b-0x00000c88,1]}", -- 0x00000c88
    x"{code[0x00000c8f-0x00000c8c,1]}", -- 0x00000c8c
    x"{code[0x00000c93-0x00000c90,1]}", -- 0x00000c90
    x"{code[0x00000c97-0x00000c94,1]}", -- 0x00000c94
    x"{code[0x00000c9b-0x00000c98,1]}", -- 0x00000c98
    x"{code[0x00000c9f-0x00000c9c,1]}", -- 0x00000c9c
    x"{code[0x00000ca3-0x00000ca0,1]}", -- 0x00000ca0
    x"{code[0x00000ca7-0x00000ca4,1]}", -- 0x00000ca4
    x"{code[0x00000cab-0x00000ca8,1]}", -- 0x00000ca8
    x"{code[0x00000caf-0x00000cac,1]}", -- 0x00000cac
    x"{code[0x00000cb3-0x00000cb0,1]}", -- 0x00000cb0
    x"{code[0x00000cb7-0x00000cb4,1]}", -- 0x00000cb4
    x"{code[0x00000cbb-0x00000cb8,1]}", -- 0x00000cb8
    x"{code[0x00000cbf-0x00000cbc,1]}", -- 0x00000cbc
    x"{code[0x00000cc3-0x00000cc0,1]}", -- 0x00000cc0
    x"{code[0x00000cc7-0x00000cc4,1]}", -- 0x00000cc4
    x"{code[0x00000ccb-0x00000cc8,1]}", -- 0x00000cc8
    x"{code[0x00000ccf-0x00000ccc,1]}", -- 0x00000ccc
    x"{code[0x00000cd3-0x00000cd0,1]}", -- 0x00000cd0
    x"{code[0x00000cd7-0x00000cd4,1]}", -- 0x00000cd4
    x"{code[0x00000cdb-0x00000cd8,1]}", -- 0x00000cd8
    x"{code[0x00000cdf-0x00000cdc,1]}", -- 0x00000cdc
    x"{code[0x00000ce3-0x00000ce0,1]}", -- 0x00000ce0
    x"{code[0x00000ce7-0x00000ce4,1]}", -- 0x00000ce4
    x"{code[0x00000ceb-0x00000ce8,1]}", -- 0x00000ce8
    x"{code[0x00000cef-0x00000cec,1]}", -- 0x00000cec
    x"{code[0x00000cf3-0x00000cf0,1]}", -- 0x00000cf0
    x"{code[0x00000cf7-0x00000cf4,1]}", -- 0x00000cf4
    x"{code[0x00000cfb-0x00000cf8,1]}", -- 0x00000cf8
    x"{code[0x00000cff-0x00000cfc,1]}", -- 0x00000cfc
    x"{code[0x00000d03-0x00000d00,1]}", -- 0x00000d00
    x"{code[0x00000d07-0x00000d04,1]}", -- 0x00000d04
    x"{code[0x00000d0b-0x00000d08,1]}", -- 0x00000d08
    x"{code[0x00000d0f-0x00000d0c,1]}", -- 0x00000d0c
    x"{code[0x00000d13-0x00000d10,1]}", -- 0x00000d10
    x"{code[0x00000d17-0x00000d14,1]}", -- 0x00000d14
    x"{code[0x00000d1b-0x00000d18,1]}", -- 0x00000d18
    x"{code[0x00000d1f-0x00000d1c,1]}", -- 0x00000d1c
    x"{code[0x00000d23-0x00000d20,1]}", -- 0x00000d20
    x"{code[0x00000d27-0x00000d24,1]}", -- 0x00000d24
    x"{code[0x00000d2b-0x00000d28,1]}", -- 0x00000d28
    x"{code[0x00000d2f-0x00000d2c,1]}", -- 0x00000d2c
    x"{code[0x00000d33-0x00000d30,1]}", -- 0x00000d30
    x"{code[0x00000d37-0x00000d34,1]}", -- 0x00000d34
    x"{code[0x00000d3b-0x00000d38,1]}", -- 0x00000d38
    x"{code[0x00000d3f-0x00000d3c,1]}", -- 0x00000d3c
    x"{code[0x00000d43-0x00000d40,1]}", -- 0x00000d40
    x"{code[0x00000d47-0x00000d44,1]}", -- 0x00000d44
    x"{code[0x00000d4b-0x00000d48,1]}", -- 0x00000d48
    x"{code[0x00000d4f-0x00000d4c,1]}", -- 0x00000d4c
    x"{code[0x00000d53-0x00000d50,1]}", -- 0x00000d50
    x"{code[0x00000d57-0x00000d54,1]}", -- 0x00000d54
    x"{code[0x00000d5b-0x00000d58,1]}", -- 0x00000d58
    x"{code[0x00000d5f-0x00000d5c,1]}", -- 0x00000d5c
    x"{code[0x00000d63-0x00000d60,1]}", -- 0x00000d60
    x"{code[0x00000d67-0x00000d64,1]}", -- 0x00000d64
    x"{code[0x00000d6b-0x00000d68,1]}", -- 0x00000d68
    x"{code[0x00000d6f-0x00000d6c,1]}", -- 0x00000d6c
    x"{code[0x00000d73-0x00000d70,1]}", -- 0x00000d70
    x"{code[0x00000d77-0x00000d74,1]}", -- 0x00000d74
    x"{code[0x00000d7b-0x00000d78,1]}", -- 0x00000d78
    x"{code[0x00000d7f-0x00000d7c,1]}", -- 0x00000d7c
    x"{code[0x00000d83-0x00000d80,1]}", -- 0x00000d80
    x"{code[0x00000d87-0x00000d84,1]}", -- 0x00000d84
    x"{code[0x00000d8b-0x00000d88,1]}", -- 0x00000d88
    x"{code[0x00000d8f-0x00000d8c,1]}", -- 0x00000d8c
    x"{code[0x00000d93-0x00000d90,1]}", -- 0x00000d90
    x"{code[0x00000d97-0x00000d94,1]}", -- 0x00000d94
    x"{code[0x00000d9b-0x00000d98,1]}", -- 0x00000d98
    x"{code[0x00000d9f-0x00000d9c,1]}", -- 0x00000d9c
    x"{code[0x00000da3-0x00000da0,1]}", -- 0x00000da0
    x"{code[0x00000da7-0x00000da4,1]}", -- 0x00000da4
    x"{code[0x00000dab-0x00000da8,1]}", -- 0x00000da8
    x"{code[0x00000daf-0x00000dac,1]}", -- 0x00000dac
    x"{code[0x00000db3-0x00000db0,1]}", -- 0x00000db0
    x"{code[0x00000db7-0x00000db4,1]}", -- 0x00000db4
    x"{code[0x00000dbb-0x00000db8,1]}", -- 0x00000db8
    x"{code[0x00000dbf-0x00000dbc,1]}", -- 0x00000dbc
    x"{code[0x00000dc3-0x00000dc0,1]}", -- 0x00000dc0
    x"{code[0x00000dc7-0x00000dc4,1]}", -- 0x00000dc4
    x"{code[0x00000dcb-0x00000dc8,1]}", -- 0x00000dc8
    x"{code[0x00000dcf-0x00000dcc,1]}", -- 0x00000dcc
    x"{code[0x00000dd3-0x00000dd0,1]}", -- 0x00000dd0
    x"{code[0x00000dd7-0x00000dd4,1]}", -- 0x00000dd4
    x"{code[0x00000ddb-0x00000dd8,1]}", -- 0x00000dd8
    x"{code[0x00000ddf-0x00000ddc,1]}", -- 0x00000ddc
    x"{code[0x00000de3-0x00000de0,1]}", -- 0x00000de0
    x"{code[0x00000de7-0x00000de4,1]}", -- 0x00000de4
    x"{code[0x00000deb-0x00000de8,1]}", -- 0x00000de8
    x"{code[0x00000def-0x00000dec,1]}", -- 0x00000dec
    x"{code[0x00000df3-0x00000df0,1]}", -- 0x00000df0
    x"{code[0x00000df7-0x00000df4,1]}", -- 0x00000df4
    x"{code[0x00000dfb-0x00000df8,1]}", -- 0x00000df8
    x"{code[0x00000dff-0x00000dfc,1]}", -- 0x00000dfc
    x"{code[0x00000e03-0x00000e00,1]}", -- 0x00000e00
    x"{code[0x00000e07-0x00000e04,1]}", -- 0x00000e04
    x"{code[0x00000e0b-0x00000e08,1]}", -- 0x00000e08
    x"{code[0x00000e0f-0x00000e0c,1]}", -- 0x00000e0c
    x"{code[0x00000e13-0x00000e10,1]}", -- 0x00000e10
    x"{code[0x00000e17-0x00000e14,1]}", -- 0x00000e14
    x"{code[0x00000e1b-0x00000e18,1]}", -- 0x00000e18
    x"{code[0x00000e1f-0x00000e1c,1]}", -- 0x00000e1c
    x"{code[0x00000e23-0x00000e20,1]}", -- 0x00000e20
    x"{code[0x00000e27-0x00000e24,1]}", -- 0x00000e24
    x"{code[0x00000e2b-0x00000e28,1]}", -- 0x00000e28
    x"{code[0x00000e2f-0x00000e2c,1]}", -- 0x00000e2c
    x"{code[0x00000e33-0x00000e30,1]}", -- 0x00000e30
    x"{code[0x00000e37-0x00000e34,1]}", -- 0x00000e34
    x"{code[0x00000e3b-0x00000e38,1]}", -- 0x00000e38
    x"{code[0x00000e3f-0x00000e3c,1]}", -- 0x00000e3c
    x"{code[0x00000e43-0x00000e40,1]}", -- 0x00000e40
    x"{code[0x00000e47-0x00000e44,1]}", -- 0x00000e44
    x"{code[0x00000e4b-0x00000e48,1]}", -- 0x00000e48
    x"{code[0x00000e4f-0x00000e4c,1]}", -- 0x00000e4c
    x"{code[0x00000e53-0x00000e50,1]}", -- 0x00000e50
    x"{code[0x00000e57-0x00000e54,1]}", -- 0x00000e54
    x"{code[0x00000e5b-0x00000e58,1]}", -- 0x00000e58
    x"{code[0x00000e5f-0x00000e5c,1]}", -- 0x00000e5c
    x"{code[0x00000e63-0x00000e60,1]}", -- 0x00000e60
    x"{code[0x00000e67-0x00000e64,1]}", -- 0x00000e64
    x"{code[0x00000e6b-0x00000e68,1]}", -- 0x00000e68
    x"{code[0x00000e6f-0x00000e6c,1]}", -- 0x00000e6c
    x"{code[0x00000e73-0x00000e70,1]}", -- 0x00000e70
    x"{code[0x00000e77-0x00000e74,1]}", -- 0x00000e74
    x"{code[0x00000e7b-0x00000e78,1]}", -- 0x00000e78
    x"{code[0x00000e7f-0x00000e7c,1]}", -- 0x00000e7c
    x"{code[0x00000e83-0x00000e80,1]}", -- 0x00000e80
    x"{code[0x00000e87-0x00000e84,1]}", -- 0x00000e84
    x"{code[0x00000e8b-0x00000e88,1]}", -- 0x00000e88
    x"{code[0x00000e8f-0x00000e8c,1]}", -- 0x00000e8c
    x"{code[0x00000e93-0x00000e90,1]}", -- 0x00000e90
    x"{code[0x00000e97-0x00000e94,1]}", -- 0x00000e94
    x"{code[0x00000e9b-0x00000e98,1]}", -- 0x00000e98
    x"{code[0x00000e9f-0x00000e9c,1]}", -- 0x00000e9c
    x"{code[0x00000ea3-0x00000ea0,1]}", -- 0x00000ea0
    x"{code[0x00000ea7-0x00000ea4,1]}", -- 0x00000ea4
    x"{code[0x00000eab-0x00000ea8,1]}", -- 0x00000ea8
    x"{code[0x00000eaf-0x00000eac,1]}", -- 0x00000eac
    x"{code[0x00000eb3-0x00000eb0,1]}", -- 0x00000eb0
    x"{code[0x00000eb7-0x00000eb4,1]}", -- 0x00000eb4
    x"{code[0x00000ebb-0x00000eb8,1]}", -- 0x00000eb8
    x"{code[0x00000ebf-0x00000ebc,1]}", -- 0x00000ebc
    x"{code[0x00000ec3-0x00000ec0,1]}", -- 0x00000ec0
    x"{code[0x00000ec7-0x00000ec4,1]}", -- 0x00000ec4
    x"{code[0x00000ecb-0x00000ec8,1]}", -- 0x00000ec8
    x"{code[0x00000ecf-0x00000ecc,1]}", -- 0x00000ecc
    x"{code[0x00000ed3-0x00000ed0,1]}", -- 0x00000ed0
    x"{code[0x00000ed7-0x00000ed4,1]}", -- 0x00000ed4
    x"{code[0x00000edb-0x00000ed8,1]}", -- 0x00000ed8
    x"{code[0x00000edf-0x00000edc,1]}", -- 0x00000edc
    x"{code[0x00000ee3-0x00000ee0,1]}", -- 0x00000ee0
    x"{code[0x00000ee7-0x00000ee4,1]}", -- 0x00000ee4
    x"{code[0x00000eeb-0x00000ee8,1]}", -- 0x00000ee8
    x"{code[0x00000eef-0x00000eec,1]}", -- 0x00000eec
    x"{code[0x00000ef3-0x00000ef0,1]}", -- 0x00000ef0
    x"{code[0x00000ef7-0x00000ef4,1]}", -- 0x00000ef4
    x"{code[0x00000efb-0x00000ef8,1]}", -- 0x00000ef8
    x"{code[0x00000eff-0x00000efc,1]}", -- 0x00000efc
    x"{code[0x00000f03-0x00000f00,1]}", -- 0x00000f00
    x"{code[0x00000f07-0x00000f04,1]}", -- 0x00000f04
    x"{code[0x00000f0b-0x00000f08,1]}", -- 0x00000f08
    x"{code[0x00000f0f-0x00000f0c,1]}", -- 0x00000f0c
    x"{code[0x00000f13-0x00000f10,1]}", -- 0x00000f10
    x"{code[0x00000f17-0x00000f14,1]}", -- 0x00000f14
    x"{code[0x00000f1b-0x00000f18,1]}", -- 0x00000f18
    x"{code[0x00000f1f-0x00000f1c,1]}", -- 0x00000f1c
    x"{code[0x00000f23-0x00000f20,1]}", -- 0x00000f20
    x"{code[0x00000f27-0x00000f24,1]}", -- 0x00000f24
    x"{code[0x00000f2b-0x00000f28,1]}", -- 0x00000f28
    x"{code[0x00000f2f-0x00000f2c,1]}", -- 0x00000f2c
    x"{code[0x00000f33-0x00000f30,1]}", -- 0x00000f30
    x"{code[0x00000f37-0x00000f34,1]}", -- 0x00000f34
    x"{code[0x00000f3b-0x00000f38,1]}", -- 0x00000f38
    x"{code[0x00000f3f-0x00000f3c,1]}", -- 0x00000f3c
    x"{code[0x00000f43-0x00000f40,1]}", -- 0x00000f40
    x"{code[0x00000f47-0x00000f44,1]}", -- 0x00000f44
    x"{code[0x00000f4b-0x00000f48,1]}", -- 0x00000f48
    x"{code[0x00000f4f-0x00000f4c,1]}", -- 0x00000f4c
    x"{code[0x00000f53-0x00000f50,1]}", -- 0x00000f50
    x"{code[0x00000f57-0x00000f54,1]}", -- 0x00000f54
    x"{code[0x00000f5b-0x00000f58,1]}", -- 0x00000f58
    x"{code[0x00000f5f-0x00000f5c,1]}", -- 0x00000f5c
    x"{code[0x00000f63-0x00000f60,1]}", -- 0x00000f60
    x"{code[0x00000f67-0x00000f64,1]}", -- 0x00000f64
    x"{code[0x00000f6b-0x00000f68,1]}", -- 0x00000f68
    x"{code[0x00000f6f-0x00000f6c,1]}", -- 0x00000f6c
    x"{code[0x00000f73-0x00000f70,1]}", -- 0x00000f70
    x"{code[0x00000f77-0x00000f74,1]}", -- 0x00000f74
    x"{code[0x00000f7b-0x00000f78,1]}", -- 0x00000f78
    x"{code[0x00000f7f-0x00000f7c,1]}", -- 0x00000f7c
    x"{code[0x00000f83-0x00000f80,1]}", -- 0x00000f80
    x"{code[0x00000f87-0x00000f84,1]}", -- 0x00000f84
    x"{code[0x00000f8b-0x00000f88,1]}", -- 0x00000f88
    x"{code[0x00000f8f-0x00000f8c,1]}", -- 0x00000f8c
    x"{code[0x00000f93-0x00000f90,1]}", -- 0x00000f90
    x"{code[0x00000f97-0x00000f94,1]}", -- 0x00000f94
    x"{code[0x00000f9b-0x00000f98,1]}", -- 0x00000f98
    x"{code[0x00000f9f-0x00000f9c,1]}", -- 0x00000f9c
    x"{code[0x00000fa3-0x00000fa0,1]}", -- 0x00000fa0
    x"{code[0x00000fa7-0x00000fa4,1]}", -- 0x00000fa4
    x"{code[0x00000fab-0x00000fa8,1]}", -- 0x00000fa8
    x"{code[0x00000faf-0x00000fac,1]}", -- 0x00000fac
    x"{code[0x00000fb3-0x00000fb0,1]}", -- 0x00000fb0
    x"{code[0x00000fb7-0x00000fb4,1]}", -- 0x00000fb4
    x"{code[0x00000fbb-0x00000fb8,1]}", -- 0x00000fb8
    x"{code[0x00000fbf-0x00000fbc,1]}", -- 0x00000fbc
    x"{code[0x00000fc3-0x00000fc0,1]}", -- 0x00000fc0
    x"{code[0x00000fc7-0x00000fc4,1]}", -- 0x00000fc4
    x"{code[0x00000fcb-0x00000fc8,1]}", -- 0x00000fc8
    x"{code[0x00000fcf-0x00000fcc,1]}", -- 0x00000fcc
    x"{code[0x00000fd3-0x00000fd0,1]}", -- 0x00000fd0
    x"{code[0x00000fd7-0x00000fd4,1]}", -- 0x00000fd4
    x"{code[0x00000fdb-0x00000fd8,1]}", -- 0x00000fd8
    x"{code[0x00000fdf-0x00000fdc,1]}", -- 0x00000fdc
    x"{code[0x00000fe3-0x00000fe0,1]}", -- 0x00000fe0
    x"{code[0x00000fe7-0x00000fe4,1]}", -- 0x00000fe4
    x"{code[0x00000feb-0x00000fe8,1]}", -- 0x00000fe8
    x"{code[0x00000fef-0x00000fec,1]}", -- 0x00000fec
    x"{code[0x00000ff3-0x00000ff0,1]}", -- 0x00000ff0
    x"{code[0x00000ff7-0x00000ff4,1]}", -- 0x00000ff4
    x"{code[0x00000ffb-0x00000ff8,1]}", -- 0x00000ff8
    x"{code[0x00000fff-0x00000ffc,1]}", -- 0x00000ffc
    x"{code[0x00001003-0x00001000,1]}", -- 0x00001000
    x"{code[0x00001007-0x00001004,1]}", -- 0x00001004
    x"{code[0x0000100b-0x00001008,1]}", -- 0x00001008
    x"{code[0x0000100f-0x0000100c,1]}", -- 0x0000100c
    x"{code[0x00001013-0x00001010,1]}", -- 0x00001010
    x"{code[0x00001017-0x00001014,1]}", -- 0x00001014
    x"{code[0x0000101b-0x00001018,1]}", -- 0x00001018
    x"{code[0x0000101f-0x0000101c,1]}", -- 0x0000101c
    x"{code[0x00001023-0x00001020,1]}", -- 0x00001020
    x"{code[0x00001027-0x00001024,1]}", -- 0x00001024
    x"{code[0x0000102b-0x00001028,1]}", -- 0x00001028
    x"{code[0x0000102f-0x0000102c,1]}", -- 0x0000102c
    x"{code[0x00001033-0x00001030,1]}", -- 0x00001030
    x"{code[0x00001037-0x00001034,1]}", -- 0x00001034
    x"{code[0x0000103b-0x00001038,1]}", -- 0x00001038
    x"{code[0x0000103f-0x0000103c,1]}", -- 0x0000103c
    x"{code[0x00001043-0x00001040,1]}", -- 0x00001040
    x"{code[0x00001047-0x00001044,1]}", -- 0x00001044
    x"{code[0x0000104b-0x00001048,1]}", -- 0x00001048
    x"{code[0x0000104f-0x0000104c,1]}", -- 0x0000104c
    x"{code[0x00001053-0x00001050,1]}", -- 0x00001050
    x"{code[0x00001057-0x00001054,1]}", -- 0x00001054
    x"{code[0x0000105b-0x00001058,1]}", -- 0x00001058
    x"{code[0x0000105f-0x0000105c,1]}", -- 0x0000105c
    x"{code[0x00001063-0x00001060,1]}", -- 0x00001060
    x"{code[0x00001067-0x00001064,1]}", -- 0x00001064
    x"{code[0x0000106b-0x00001068,1]}", -- 0x00001068
    x"{code[0x0000106f-0x0000106c,1]}", -- 0x0000106c
    x"{code[0x00001073-0x00001070,1]}", -- 0x00001070
    x"{code[0x00001077-0x00001074,1]}", -- 0x00001074
    x"{code[0x0000107b-0x00001078,1]}", -- 0x00001078
    x"{code[0x0000107f-0x0000107c,1]}", -- 0x0000107c
    x"{code[0x00001083-0x00001080,1]}", -- 0x00001080
    x"{code[0x00001087-0x00001084,1]}", -- 0x00001084
    x"{code[0x0000108b-0x00001088,1]}", -- 0x00001088
    x"{code[0x0000108f-0x0000108c,1]}", -- 0x0000108c
    x"{code[0x00001093-0x00001090,1]}", -- 0x00001090
    x"{code[0x00001097-0x00001094,1]}", -- 0x00001094
    x"{code[0x0000109b-0x00001098,1]}", -- 0x00001098
    x"{code[0x0000109f-0x0000109c,1]}", -- 0x0000109c
    x"{code[0x000010a3-0x000010a0,1]}", -- 0x000010a0
    x"{code[0x000010a7-0x000010a4,1]}", -- 0x000010a4
    x"{code[0x000010ab-0x000010a8,1]}", -- 0x000010a8
    x"{code[0x000010af-0x000010ac,1]}", -- 0x000010ac
    x"{code[0x000010b3-0x000010b0,1]}", -- 0x000010b0
    x"{code[0x000010b7-0x000010b4,1]}", -- 0x000010b4
    x"{code[0x000010bb-0x000010b8,1]}", -- 0x000010b8
    x"{code[0x000010bf-0x000010bc,1]}", -- 0x000010bc
    x"{code[0x000010c3-0x000010c0,1]}", -- 0x000010c0
    x"{code[0x000010c7-0x000010c4,1]}", -- 0x000010c4
    x"{code[0x000010cb-0x000010c8,1]}", -- 0x000010c8
    x"{code[0x000010cf-0x000010cc,1]}", -- 0x000010cc
    x"{code[0x000010d3-0x000010d0,1]}", -- 0x000010d0
    x"{code[0x000010d7-0x000010d4,1]}", -- 0x000010d4
    x"{code[0x000010db-0x000010d8,1]}", -- 0x000010d8
    x"{code[0x000010df-0x000010dc,1]}", -- 0x000010dc
    x"{code[0x000010e3-0x000010e0,1]}", -- 0x000010e0
    x"{code[0x000010e7-0x000010e4,1]}", -- 0x000010e4
    x"{code[0x000010eb-0x000010e8,1]}", -- 0x000010e8
    x"{code[0x000010ef-0x000010ec,1]}", -- 0x000010ec
    x"{code[0x000010f3-0x000010f0,1]}", -- 0x000010f0
    x"{code[0x000010f7-0x000010f4,1]}", -- 0x000010f4
    x"{code[0x000010fb-0x000010f8,1]}", -- 0x000010f8
    x"{code[0x000010ff-0x000010fc,1]}", -- 0x000010fc
    x"{code[0x00001103-0x00001100,1]}", -- 0x00001100
    x"{code[0x00001107-0x00001104,1]}", -- 0x00001104
    x"{code[0x0000110b-0x00001108,1]}", -- 0x00001108
    x"{code[0x0000110f-0x0000110c,1]}", -- 0x0000110c
    x"{code[0x00001113-0x00001110,1]}", -- 0x00001110
    x"{code[0x00001117-0x00001114,1]}", -- 0x00001114
    x"{code[0x0000111b-0x00001118,1]}", -- 0x00001118
    x"{code[0x0000111f-0x0000111c,1]}", -- 0x0000111c
    x"{code[0x00001123-0x00001120,1]}", -- 0x00001120
    x"{code[0x00001127-0x00001124,1]}", -- 0x00001124
    x"{code[0x0000112b-0x00001128,1]}", -- 0x00001128
    x"{code[0x0000112f-0x0000112c,1]}", -- 0x0000112c
    x"{code[0x00001133-0x00001130,1]}", -- 0x00001130
    x"{code[0x00001137-0x00001134,1]}", -- 0x00001134
    x"{code[0x0000113b-0x00001138,1]}", -- 0x00001138
    x"{code[0x0000113f-0x0000113c,1]}", -- 0x0000113c
    x"{code[0x00001143-0x00001140,1]}", -- 0x00001140
    x"{code[0x00001147-0x00001144,1]}", -- 0x00001144
    x"{code[0x0000114b-0x00001148,1]}", -- 0x00001148
    x"{code[0x0000114f-0x0000114c,1]}", -- 0x0000114c
    x"{code[0x00001153-0x00001150,1]}", -- 0x00001150
    x"{code[0x00001157-0x00001154,1]}", -- 0x00001154
    x"{code[0x0000115b-0x00001158,1]}", -- 0x00001158
    x"{code[0x0000115f-0x0000115c,1]}", -- 0x0000115c
    x"{code[0x00001163-0x00001160,1]}", -- 0x00001160
    x"{code[0x00001167-0x00001164,1]}", -- 0x00001164
    x"{code[0x0000116b-0x00001168,1]}", -- 0x00001168
    x"{code[0x0000116f-0x0000116c,1]}", -- 0x0000116c
    x"{code[0x00001173-0x00001170,1]}", -- 0x00001170
    x"{code[0x00001177-0x00001174,1]}", -- 0x00001174
    x"{code[0x0000117b-0x00001178,1]}", -- 0x00001178
    x"{code[0x0000117f-0x0000117c,1]}", -- 0x0000117c
    x"{code[0x00001183-0x00001180,1]}", -- 0x00001180
    x"{code[0x00001187-0x00001184,1]}", -- 0x00001184
    x"{code[0x0000118b-0x00001188,1]}", -- 0x00001188
    x"{code[0x0000118f-0x0000118c,1]}", -- 0x0000118c
    x"{code[0x00001193-0x00001190,1]}", -- 0x00001190
    x"{code[0x00001197-0x00001194,1]}", -- 0x00001194
    x"{code[0x0000119b-0x00001198,1]}", -- 0x00001198
    x"{code[0x0000119f-0x0000119c,1]}", -- 0x0000119c
    x"{code[0x000011a3-0x000011a0,1]}", -- 0x000011a0
    x"{code[0x000011a7-0x000011a4,1]}", -- 0x000011a4
    x"{code[0x000011ab-0x000011a8,1]}", -- 0x000011a8
    x"{code[0x000011af-0x000011ac,1]}", -- 0x000011ac
    x"{code[0x000011b3-0x000011b0,1]}", -- 0x000011b0
    x"{code[0x000011b7-0x000011b4,1]}", -- 0x000011b4
    x"{code[0x000011bb-0x000011b8,1]}", -- 0x000011b8
    x"{code[0x000011bf-0x000011bc,1]}", -- 0x000011bc
    x"{code[0x000011c3-0x000011c0,1]}", -- 0x000011c0
    x"{code[0x000011c7-0x000011c4,1]}", -- 0x000011c4
    x"{code[0x000011cb-0x000011c8,1]}", -- 0x000011c8
    x"{code[0x000011cf-0x000011cc,1]}", -- 0x000011cc
    x"{code[0x000011d3-0x000011d0,1]}", -- 0x000011d0
    x"{code[0x000011d7-0x000011d4,1]}", -- 0x000011d4
    x"{code[0x000011db-0x000011d8,1]}", -- 0x000011d8
    x"{code[0x000011df-0x000011dc,1]}", -- 0x000011dc
    x"{code[0x000011e3-0x000011e0,1]}", -- 0x000011e0
    x"{code[0x000011e7-0x000011e4,1]}", -- 0x000011e4
    x"{code[0x000011eb-0x000011e8,1]}", -- 0x000011e8
    x"{code[0x000011ef-0x000011ec,1]}", -- 0x000011ec
    x"{code[0x000011f3-0x000011f0,1]}", -- 0x000011f0
    x"{code[0x000011f7-0x000011f4,1]}", -- 0x000011f4
    x"{code[0x000011fb-0x000011f8,1]}", -- 0x000011f8
    x"{code[0x000011ff-0x000011fc,1]}", -- 0x000011fc
    x"{code[0x00001203-0x00001200,1]}", -- 0x00001200
    x"{code[0x00001207-0x00001204,1]}", -- 0x00001204
    x"{code[0x0000120b-0x00001208,1]}", -- 0x00001208
    x"{code[0x0000120f-0x0000120c,1]}", -- 0x0000120c
    x"{code[0x00001213-0x00001210,1]}", -- 0x00001210
    x"{code[0x00001217-0x00001214,1]}", -- 0x00001214
    x"{code[0x0000121b-0x00001218,1]}", -- 0x00001218
    x"{code[0x0000121f-0x0000121c,1]}", -- 0x0000121c
    x"{code[0x00001223-0x00001220,1]}", -- 0x00001220
    x"{code[0x00001227-0x00001224,1]}", -- 0x00001224
    x"{code[0x0000122b-0x00001228,1]}", -- 0x00001228
    x"{code[0x0000122f-0x0000122c,1]}", -- 0x0000122c
    x"{code[0x00001233-0x00001230,1]}", -- 0x00001230
    x"{code[0x00001237-0x00001234,1]}", -- 0x00001234
    x"{code[0x0000123b-0x00001238,1]}", -- 0x00001238
    x"{code[0x0000123f-0x0000123c,1]}", -- 0x0000123c
    x"{code[0x00001243-0x00001240,1]}", -- 0x00001240
    x"{code[0x00001247-0x00001244,1]}", -- 0x00001244
    x"{code[0x0000124b-0x00001248,1]}", -- 0x00001248
    x"{code[0x0000124f-0x0000124c,1]}", -- 0x0000124c
    x"{code[0x00001253-0x00001250,1]}", -- 0x00001250
    x"{code[0x00001257-0x00001254,1]}", -- 0x00001254
    x"{code[0x0000125b-0x00001258,1]}", -- 0x00001258
    x"{code[0x0000125f-0x0000125c,1]}", -- 0x0000125c
    x"{code[0x00001263-0x00001260,1]}", -- 0x00001260
    x"{code[0x00001267-0x00001264,1]}", -- 0x00001264
    x"{code[0x0000126b-0x00001268,1]}", -- 0x00001268
    x"{code[0x0000126f-0x0000126c,1]}", -- 0x0000126c
    x"{code[0x00001273-0x00001270,1]}", -- 0x00001270
    x"{code[0x00001277-0x00001274,1]}", -- 0x00001274
    x"{code[0x0000127b-0x00001278,1]}", -- 0x00001278
    x"{code[0x0000127f-0x0000127c,1]}", -- 0x0000127c
    x"{code[0x00001283-0x00001280,1]}", -- 0x00001280
    x"{code[0x00001287-0x00001284,1]}", -- 0x00001284
    x"{code[0x0000128b-0x00001288,1]}", -- 0x00001288
    x"{code[0x0000128f-0x0000128c,1]}", -- 0x0000128c
    x"{code[0x00001293-0x00001290,1]}", -- 0x00001290
    x"{code[0x00001297-0x00001294,1]}", -- 0x00001294
    x"{code[0x0000129b-0x00001298,1]}", -- 0x00001298
    x"{code[0x0000129f-0x0000129c,1]}", -- 0x0000129c
    x"{code[0x000012a3-0x000012a0,1]}", -- 0x000012a0
    x"{code[0x000012a7-0x000012a4,1]}", -- 0x000012a4
    x"{code[0x000012ab-0x000012a8,1]}", -- 0x000012a8
    x"{code[0x000012af-0x000012ac,1]}", -- 0x000012ac
    x"{code[0x000012b3-0x000012b0,1]}", -- 0x000012b0
    x"{code[0x000012b7-0x000012b4,1]}", -- 0x000012b4
    x"{code[0x000012bb-0x000012b8,1]}", -- 0x000012b8
    x"{code[0x000012bf-0x000012bc,1]}", -- 0x000012bc
    x"{code[0x000012c3-0x000012c0,1]}", -- 0x000012c0
    x"{code[0x000012c7-0x000012c4,1]}", -- 0x000012c4
    x"{code[0x000012cb-0x000012c8,1]}", -- 0x000012c8
    x"{code[0x000012cf-0x000012cc,1]}", -- 0x000012cc
    x"{code[0x000012d3-0x000012d0,1]}", -- 0x000012d0
    x"{code[0x000012d7-0x000012d4,1]}", -- 0x000012d4
    x"{code[0x000012db-0x000012d8,1]}", -- 0x000012d8
    x"{code[0x000012df-0x000012dc,1]}", -- 0x000012dc
    x"{code[0x000012e3-0x000012e0,1]}", -- 0x000012e0
    x"{code[0x000012e7-0x000012e4,1]}", -- 0x000012e4
    x"{code[0x000012eb-0x000012e8,1]}", -- 0x000012e8
    x"{code[0x000012ef-0x000012ec,1]}", -- 0x000012ec
    x"{code[0x000012f3-0x000012f0,1]}", -- 0x000012f0
    x"{code[0x000012f7-0x000012f4,1]}", -- 0x000012f4
    x"{code[0x000012fb-0x000012f8,1]}", -- 0x000012f8
    x"{code[0x000012ff-0x000012fc,1]}", -- 0x000012fc
    x"{code[0x00001303-0x00001300,1]}", -- 0x00001300
    x"{code[0x00001307-0x00001304,1]}", -- 0x00001304
    x"{code[0x0000130b-0x00001308,1]}", -- 0x00001308
    x"{code[0x0000130f-0x0000130c,1]}", -- 0x0000130c
    x"{code[0x00001313-0x00001310,1]}", -- 0x00001310
    x"{code[0x00001317-0x00001314,1]}", -- 0x00001314
    x"{code[0x0000131b-0x00001318,1]}", -- 0x00001318
    x"{code[0x0000131f-0x0000131c,1]}", -- 0x0000131c
    x"{code[0x00001323-0x00001320,1]}", -- 0x00001320
    x"{code[0x00001327-0x00001324,1]}", -- 0x00001324
    x"{code[0x0000132b-0x00001328,1]}", -- 0x00001328
    x"{code[0x0000132f-0x0000132c,1]}", -- 0x0000132c
    x"{code[0x00001333-0x00001330,1]}", -- 0x00001330
    x"{code[0x00001337-0x00001334,1]}", -- 0x00001334
    x"{code[0x0000133b-0x00001338,1]}", -- 0x00001338
    x"{code[0x0000133f-0x0000133c,1]}", -- 0x0000133c
    x"{code[0x00001343-0x00001340,1]}", -- 0x00001340
    x"{code[0x00001347-0x00001344,1]}", -- 0x00001344
    x"{code[0x0000134b-0x00001348,1]}", -- 0x00001348
    x"{code[0x0000134f-0x0000134c,1]}", -- 0x0000134c
    x"{code[0x00001353-0x00001350,1]}", -- 0x00001350
    x"{code[0x00001357-0x00001354,1]}", -- 0x00001354
    x"{code[0x0000135b-0x00001358,1]}", -- 0x00001358
    x"{code[0x0000135f-0x0000135c,1]}", -- 0x0000135c
    x"{code[0x00001363-0x00001360,1]}", -- 0x00001360
    x"{code[0x00001367-0x00001364,1]}", -- 0x00001364
    x"{code[0x0000136b-0x00001368,1]}", -- 0x00001368
    x"{code[0x0000136f-0x0000136c,1]}", -- 0x0000136c
    x"{code[0x00001373-0x00001370,1]}", -- 0x00001370
    x"{code[0x00001377-0x00001374,1]}", -- 0x00001374
    x"{code[0x0000137b-0x00001378,1]}", -- 0x00001378
    x"{code[0x0000137f-0x0000137c,1]}", -- 0x0000137c
    x"{code[0x00001383-0x00001380,1]}", -- 0x00001380
    x"{code[0x00001387-0x00001384,1]}", -- 0x00001384
    x"{code[0x0000138b-0x00001388,1]}", -- 0x00001388
    x"{code[0x0000138f-0x0000138c,1]}", -- 0x0000138c
    x"{code[0x00001393-0x00001390,1]}", -- 0x00001390
    x"{code[0x00001397-0x00001394,1]}", -- 0x00001394
    x"{code[0x0000139b-0x00001398,1]}", -- 0x00001398
    x"{code[0x0000139f-0x0000139c,1]}", -- 0x0000139c
    x"{code[0x000013a3-0x000013a0,1]}", -- 0x000013a0
    x"{code[0x000013a7-0x000013a4,1]}", -- 0x000013a4
    x"{code[0x000013ab-0x000013a8,1]}", -- 0x000013a8
    x"{code[0x000013af-0x000013ac,1]}", -- 0x000013ac
    x"{code[0x000013b3-0x000013b0,1]}", -- 0x000013b0
    x"{code[0x000013b7-0x000013b4,1]}", -- 0x000013b4
    x"{code[0x000013bb-0x000013b8,1]}", -- 0x000013b8
    x"{code[0x000013bf-0x000013bc,1]}", -- 0x000013bc
    x"{code[0x000013c3-0x000013c0,1]}", -- 0x000013c0
    x"{code[0x000013c7-0x000013c4,1]}", -- 0x000013c4
    x"{code[0x000013cb-0x000013c8,1]}", -- 0x000013c8
    x"{code[0x000013cf-0x000013cc,1]}", -- 0x000013cc
    x"{code[0x000013d3-0x000013d0,1]}", -- 0x000013d0
    x"{code[0x000013d7-0x000013d4,1]}", -- 0x000013d4
    x"{code[0x000013db-0x000013d8,1]}", -- 0x000013d8
    x"{code[0x000013df-0x000013dc,1]}", -- 0x000013dc
    x"{code[0x000013e3-0x000013e0,1]}", -- 0x000013e0
    x"{code[0x000013e7-0x000013e4,1]}", -- 0x000013e4
    x"{code[0x000013eb-0x000013e8,1]}", -- 0x000013e8
    x"{code[0x000013ef-0x000013ec,1]}", -- 0x000013ec
    x"{code[0x000013f3-0x000013f0,1]}", -- 0x000013f0
    x"{code[0x000013f7-0x000013f4,1]}", -- 0x000013f4
    x"{code[0x000013fb-0x000013f8,1]}", -- 0x000013f8
    x"{code[0x000013ff-0x000013fc,1]}", -- 0x000013fc
    x"{code[0x00001403-0x00001400,1]}", -- 0x00001400
    x"{code[0x00001407-0x00001404,1]}", -- 0x00001404
    x"{code[0x0000140b-0x00001408,1]}", -- 0x00001408
    x"{code[0x0000140f-0x0000140c,1]}", -- 0x0000140c
    x"{code[0x00001413-0x00001410,1]}", -- 0x00001410
    x"{code[0x00001417-0x00001414,1]}", -- 0x00001414
    x"{code[0x0000141b-0x00001418,1]}", -- 0x00001418
    x"{code[0x0000141f-0x0000141c,1]}", -- 0x0000141c
    x"{code[0x00001423-0x00001420,1]}", -- 0x00001420
    x"{code[0x00001427-0x00001424,1]}", -- 0x00001424
    x"{code[0x0000142b-0x00001428,1]}", -- 0x00001428
    x"{code[0x0000142f-0x0000142c,1]}", -- 0x0000142c
    x"{code[0x00001433-0x00001430,1]}", -- 0x00001430
    x"{code[0x00001437-0x00001434,1]}", -- 0x00001434
    x"{code[0x0000143b-0x00001438,1]}", -- 0x00001438
    x"{code[0x0000143f-0x0000143c,1]}", -- 0x0000143c
    x"{code[0x00001443-0x00001440,1]}", -- 0x00001440
    x"{code[0x00001447-0x00001444,1]}", -- 0x00001444
    x"{code[0x0000144b-0x00001448,1]}", -- 0x00001448
    x"{code[0x0000144f-0x0000144c,1]}", -- 0x0000144c
    x"{code[0x00001453-0x00001450,1]}", -- 0x00001450
    x"{code[0x00001457-0x00001454,1]}", -- 0x00001454
    x"{code[0x0000145b-0x00001458,1]}", -- 0x00001458
    x"{code[0x0000145f-0x0000145c,1]}", -- 0x0000145c
    x"{code[0x00001463-0x00001460,1]}", -- 0x00001460
    x"{code[0x00001467-0x00001464,1]}", -- 0x00001464
    x"{code[0x0000146b-0x00001468,1]}", -- 0x00001468
    x"{code[0x0000146f-0x0000146c,1]}", -- 0x0000146c
    x"{code[0x00001473-0x00001470,1]}", -- 0x00001470
    x"{code[0x00001477-0x00001474,1]}", -- 0x00001474
    x"{code[0x0000147b-0x00001478,1]}", -- 0x00001478
    x"{code[0x0000147f-0x0000147c,1]}", -- 0x0000147c
    x"{code[0x00001483-0x00001480,1]}", -- 0x00001480
    x"{code[0x00001487-0x00001484,1]}", -- 0x00001484
    x"{code[0x0000148b-0x00001488,1]}", -- 0x00001488
    x"{code[0x0000148f-0x0000148c,1]}", -- 0x0000148c
    x"{code[0x00001493-0x00001490,1]}", -- 0x00001490
    x"{code[0x00001497-0x00001494,1]}", -- 0x00001494
    x"{code[0x0000149b-0x00001498,1]}", -- 0x00001498
    x"{code[0x0000149f-0x0000149c,1]}", -- 0x0000149c
    x"{code[0x000014a3-0x000014a0,1]}", -- 0x000014a0
    x"{code[0x000014a7-0x000014a4,1]}", -- 0x000014a4
    x"{code[0x000014ab-0x000014a8,1]}", -- 0x000014a8
    x"{code[0x000014af-0x000014ac,1]}", -- 0x000014ac
    x"{code[0x000014b3-0x000014b0,1]}", -- 0x000014b0
    x"{code[0x000014b7-0x000014b4,1]}", -- 0x000014b4
    x"{code[0x000014bb-0x000014b8,1]}", -- 0x000014b8
    x"{code[0x000014bf-0x000014bc,1]}", -- 0x000014bc
    x"{code[0x000014c3-0x000014c0,1]}", -- 0x000014c0
    x"{code[0x000014c7-0x000014c4,1]}", -- 0x000014c4
    x"{code[0x000014cb-0x000014c8,1]}", -- 0x000014c8
    x"{code[0x000014cf-0x000014cc,1]}", -- 0x000014cc
    x"{code[0x000014d3-0x000014d0,1]}", -- 0x000014d0
    x"{code[0x000014d7-0x000014d4,1]}", -- 0x000014d4
    x"{code[0x000014db-0x000014d8,1]}", -- 0x000014d8
    x"{code[0x000014df-0x000014dc,1]}", -- 0x000014dc
    x"{code[0x000014e3-0x000014e0,1]}", -- 0x000014e0
    x"{code[0x000014e7-0x000014e4,1]}", -- 0x000014e4
    x"{code[0x000014eb-0x000014e8,1]}", -- 0x000014e8
    x"{code[0x000014ef-0x000014ec,1]}", -- 0x000014ec
    x"{code[0x000014f3-0x000014f0,1]}", -- 0x000014f0
    x"{code[0x000014f7-0x000014f4,1]}", -- 0x000014f4
    x"{code[0x000014fb-0x000014f8,1]}", -- 0x000014f8
    x"{code[0x000014ff-0x000014fc,1]}", -- 0x000014fc
    x"{code[0x00001503-0x00001500,1]}", -- 0x00001500
    x"{code[0x00001507-0x00001504,1]}", -- 0x00001504
    x"{code[0x0000150b-0x00001508,1]}", -- 0x00001508
    x"{code[0x0000150f-0x0000150c,1]}", -- 0x0000150c
    x"{code[0x00001513-0x00001510,1]}", -- 0x00001510
    x"{code[0x00001517-0x00001514,1]}", -- 0x00001514
    x"{code[0x0000151b-0x00001518,1]}", -- 0x00001518
    x"{code[0x0000151f-0x0000151c,1]}", -- 0x0000151c
    x"{code[0x00001523-0x00001520,1]}", -- 0x00001520
    x"{code[0x00001527-0x00001524,1]}", -- 0x00001524
    x"{code[0x0000152b-0x00001528,1]}", -- 0x00001528
    x"{code[0x0000152f-0x0000152c,1]}", -- 0x0000152c
    x"{code[0x00001533-0x00001530,1]}", -- 0x00001530
    x"{code[0x00001537-0x00001534,1]}", -- 0x00001534
    x"{code[0x0000153b-0x00001538,1]}", -- 0x00001538
    x"{code[0x0000153f-0x0000153c,1]}", -- 0x0000153c
    x"{code[0x00001543-0x00001540,1]}", -- 0x00001540
    x"{code[0x00001547-0x00001544,1]}", -- 0x00001544
    x"{code[0x0000154b-0x00001548,1]}", -- 0x00001548
    x"{code[0x0000154f-0x0000154c,1]}", -- 0x0000154c
    x"{code[0x00001553-0x00001550,1]}", -- 0x00001550
    x"{code[0x00001557-0x00001554,1]}", -- 0x00001554
    x"{code[0x0000155b-0x00001558,1]}", -- 0x00001558
    x"{code[0x0000155f-0x0000155c,1]}", -- 0x0000155c
    x"{code[0x00001563-0x00001560,1]}", -- 0x00001560
    x"{code[0x00001567-0x00001564,1]}", -- 0x00001564
    x"{code[0x0000156b-0x00001568,1]}", -- 0x00001568
    x"{code[0x0000156f-0x0000156c,1]}", -- 0x0000156c
    x"{code[0x00001573-0x00001570,1]}", -- 0x00001570
    x"{code[0x00001577-0x00001574,1]}", -- 0x00001574
    x"{code[0x0000157b-0x00001578,1]}", -- 0x00001578
    x"{code[0x0000157f-0x0000157c,1]}", -- 0x0000157c
    x"{code[0x00001583-0x00001580,1]}", -- 0x00001580
    x"{code[0x00001587-0x00001584,1]}", -- 0x00001584
    x"{code[0x0000158b-0x00001588,1]}", -- 0x00001588
    x"{code[0x0000158f-0x0000158c,1]}", -- 0x0000158c
    x"{code[0x00001593-0x00001590,1]}", -- 0x00001590
    x"{code[0x00001597-0x00001594,1]}", -- 0x00001594
    x"{code[0x0000159b-0x00001598,1]}", -- 0x00001598
    x"{code[0x0000159f-0x0000159c,1]}", -- 0x0000159c
    x"{code[0x000015a3-0x000015a0,1]}", -- 0x000015a0
    x"{code[0x000015a7-0x000015a4,1]}", -- 0x000015a4
    x"{code[0x000015ab-0x000015a8,1]}", -- 0x000015a8
    x"{code[0x000015af-0x000015ac,1]}", -- 0x000015ac
    x"{code[0x000015b3-0x000015b0,1]}", -- 0x000015b0
    x"{code[0x000015b7-0x000015b4,1]}", -- 0x000015b4
    x"{code[0x000015bb-0x000015b8,1]}", -- 0x000015b8
    x"{code[0x000015bf-0x000015bc,1]}", -- 0x000015bc
    x"{code[0x000015c3-0x000015c0,1]}", -- 0x000015c0
    x"{code[0x000015c7-0x000015c4,1]}", -- 0x000015c4
    x"{code[0x000015cb-0x000015c8,1]}", -- 0x000015c8
    x"{code[0x000015cf-0x000015cc,1]}", -- 0x000015cc
    x"{code[0x000015d3-0x000015d0,1]}", -- 0x000015d0
    x"{code[0x000015d7-0x000015d4,1]}", -- 0x000015d4
    x"{code[0x000015db-0x000015d8,1]}", -- 0x000015d8
    x"{code[0x000015df-0x000015dc,1]}", -- 0x000015dc
    x"{code[0x000015e3-0x000015e0,1]}", -- 0x000015e0
    x"{code[0x000015e7-0x000015e4,1]}", -- 0x000015e4
    x"{code[0x000015eb-0x000015e8,1]}", -- 0x000015e8
    x"{code[0x000015ef-0x000015ec,1]}", -- 0x000015ec
    x"{code[0x000015f3-0x000015f0,1]}", -- 0x000015f0
    x"{code[0x000015f7-0x000015f4,1]}", -- 0x000015f4
    x"{code[0x000015fb-0x000015f8,1]}", -- 0x000015f8
    x"{code[0x000015ff-0x000015fc,1]}", -- 0x000015fc
    x"{code[0x00001603-0x00001600,1]}", -- 0x00001600
    x"{code[0x00001607-0x00001604,1]}", -- 0x00001604
    x"{code[0x0000160b-0x00001608,1]}", -- 0x00001608
    x"{code[0x0000160f-0x0000160c,1]}", -- 0x0000160c
    x"{code[0x00001613-0x00001610,1]}", -- 0x00001610
    x"{code[0x00001617-0x00001614,1]}", -- 0x00001614
    x"{code[0x0000161b-0x00001618,1]}", -- 0x00001618
    x"{code[0x0000161f-0x0000161c,1]}", -- 0x0000161c
    x"{code[0x00001623-0x00001620,1]}", -- 0x00001620
    x"{code[0x00001627-0x00001624,1]}", -- 0x00001624
    x"{code[0x0000162b-0x00001628,1]}", -- 0x00001628
    x"{code[0x0000162f-0x0000162c,1]}", -- 0x0000162c
    x"{code[0x00001633-0x00001630,1]}", -- 0x00001630
    x"{code[0x00001637-0x00001634,1]}", -- 0x00001634
    x"{code[0x0000163b-0x00001638,1]}", -- 0x00001638
    x"{code[0x0000163f-0x0000163c,1]}", -- 0x0000163c
    x"{code[0x00001643-0x00001640,1]}", -- 0x00001640
    x"{code[0x00001647-0x00001644,1]}", -- 0x00001644
    x"{code[0x0000164b-0x00001648,1]}", -- 0x00001648
    x"{code[0x0000164f-0x0000164c,1]}", -- 0x0000164c
    x"{code[0x00001653-0x00001650,1]}", -- 0x00001650
    x"{code[0x00001657-0x00001654,1]}", -- 0x00001654
    x"{code[0x0000165b-0x00001658,1]}", -- 0x00001658
    x"{code[0x0000165f-0x0000165c,1]}", -- 0x0000165c
    x"{code[0x00001663-0x00001660,1]}", -- 0x00001660
    x"{code[0x00001667-0x00001664,1]}", -- 0x00001664
    x"{code[0x0000166b-0x00001668,1]}", -- 0x00001668
    x"{code[0x0000166f-0x0000166c,1]}", -- 0x0000166c
    x"{code[0x00001673-0x00001670,1]}", -- 0x00001670
    x"{code[0x00001677-0x00001674,1]}", -- 0x00001674
    x"{code[0x0000167b-0x00001678,1]}", -- 0x00001678
    x"{code[0x0000167f-0x0000167c,1]}", -- 0x0000167c
    x"{code[0x00001683-0x00001680,1]}", -- 0x00001680
    x"{code[0x00001687-0x00001684,1]}", -- 0x00001684
    x"{code[0x0000168b-0x00001688,1]}", -- 0x00001688
    x"{code[0x0000168f-0x0000168c,1]}", -- 0x0000168c
    x"{code[0x00001693-0x00001690,1]}", -- 0x00001690
    x"{code[0x00001697-0x00001694,1]}", -- 0x00001694
    x"{code[0x0000169b-0x00001698,1]}", -- 0x00001698
    x"{code[0x0000169f-0x0000169c,1]}", -- 0x0000169c
    x"{code[0x000016a3-0x000016a0,1]}", -- 0x000016a0
    x"{code[0x000016a7-0x000016a4,1]}", -- 0x000016a4
    x"{code[0x000016ab-0x000016a8,1]}", -- 0x000016a8
    x"{code[0x000016af-0x000016ac,1]}", -- 0x000016ac
    x"{code[0x000016b3-0x000016b0,1]}", -- 0x000016b0
    x"{code[0x000016b7-0x000016b4,1]}", -- 0x000016b4
    x"{code[0x000016bb-0x000016b8,1]}", -- 0x000016b8
    x"{code[0x000016bf-0x000016bc,1]}", -- 0x000016bc
    x"{code[0x000016c3-0x000016c0,1]}", -- 0x000016c0
    x"{code[0x000016c7-0x000016c4,1]}", -- 0x000016c4
    x"{code[0x000016cb-0x000016c8,1]}", -- 0x000016c8
    x"{code[0x000016cf-0x000016cc,1]}", -- 0x000016cc
    x"{code[0x000016d3-0x000016d0,1]}", -- 0x000016d0
    x"{code[0x000016d7-0x000016d4,1]}", -- 0x000016d4
    x"{code[0x000016db-0x000016d8,1]}", -- 0x000016d8
    x"{code[0x000016df-0x000016dc,1]}", -- 0x000016dc
    x"{code[0x000016e3-0x000016e0,1]}", -- 0x000016e0
    x"{code[0x000016e7-0x000016e4,1]}", -- 0x000016e4
    x"{code[0x000016eb-0x000016e8,1]}", -- 0x000016e8
    x"{code[0x000016ef-0x000016ec,1]}", -- 0x000016ec
    x"{code[0x000016f3-0x000016f0,1]}", -- 0x000016f0
    x"{code[0x000016f7-0x000016f4,1]}", -- 0x000016f4
    x"{code[0x000016fb-0x000016f8,1]}", -- 0x000016f8
    x"{code[0x000016ff-0x000016fc,1]}", -- 0x000016fc
    x"{code[0x00001703-0x00001700,1]}", -- 0x00001700
    x"{code[0x00001707-0x00001704,1]}", -- 0x00001704
    x"{code[0x0000170b-0x00001708,1]}", -- 0x00001708
    x"{code[0x0000170f-0x0000170c,1]}", -- 0x0000170c
    x"{code[0x00001713-0x00001710,1]}", -- 0x00001710
    x"{code[0x00001717-0x00001714,1]}", -- 0x00001714
    x"{code[0x0000171b-0x00001718,1]}", -- 0x00001718
    x"{code[0x0000171f-0x0000171c,1]}", -- 0x0000171c
    x"{code[0x00001723-0x00001720,1]}", -- 0x00001720
    x"{code[0x00001727-0x00001724,1]}", -- 0x00001724
    x"{code[0x0000172b-0x00001728,1]}", -- 0x00001728
    x"{code[0x0000172f-0x0000172c,1]}", -- 0x0000172c
    x"{code[0x00001733-0x00001730,1]}", -- 0x00001730
    x"{code[0x00001737-0x00001734,1]}", -- 0x00001734
    x"{code[0x0000173b-0x00001738,1]}", -- 0x00001738
    x"{code[0x0000173f-0x0000173c,1]}", -- 0x0000173c
    x"{code[0x00001743-0x00001740,1]}", -- 0x00001740
    x"{code[0x00001747-0x00001744,1]}", -- 0x00001744
    x"{code[0x0000174b-0x00001748,1]}", -- 0x00001748
    x"{code[0x0000174f-0x0000174c,1]}", -- 0x0000174c
    x"{code[0x00001753-0x00001750,1]}", -- 0x00001750
    x"{code[0x00001757-0x00001754,1]}", -- 0x00001754
    x"{code[0x0000175b-0x00001758,1]}", -- 0x00001758
    x"{code[0x0000175f-0x0000175c,1]}", -- 0x0000175c
    x"{code[0x00001763-0x00001760,1]}", -- 0x00001760
    x"{code[0x00001767-0x00001764,1]}", -- 0x00001764
    x"{code[0x0000176b-0x00001768,1]}", -- 0x00001768
    x"{code[0x0000176f-0x0000176c,1]}", -- 0x0000176c
    x"{code[0x00001773-0x00001770,1]}", -- 0x00001770
    x"{code[0x00001777-0x00001774,1]}", -- 0x00001774
    x"{code[0x0000177b-0x00001778,1]}", -- 0x00001778
    x"{code[0x0000177f-0x0000177c,1]}", -- 0x0000177c
    x"{code[0x00001783-0x00001780,1]}", -- 0x00001780
    x"{code[0x00001787-0x00001784,1]}", -- 0x00001784
    x"{code[0x0000178b-0x00001788,1]}", -- 0x00001788
    x"{code[0x0000178f-0x0000178c,1]}", -- 0x0000178c
    x"{code[0x00001793-0x00001790,1]}", -- 0x00001790
    x"{code[0x00001797-0x00001794,1]}", -- 0x00001794
    x"{code[0x0000179b-0x00001798,1]}", -- 0x00001798
    x"{code[0x0000179f-0x0000179c,1]}", -- 0x0000179c
    x"{code[0x000017a3-0x000017a0,1]}", -- 0x000017a0
    x"{code[0x000017a7-0x000017a4,1]}", -- 0x000017a4
    x"{code[0x000017ab-0x000017a8,1]}", -- 0x000017a8
    x"{code[0x000017af-0x000017ac,1]}", -- 0x000017ac
    x"{code[0x000017b3-0x000017b0,1]}", -- 0x000017b0
    x"{code[0x000017b7-0x000017b4,1]}", -- 0x000017b4
    x"{code[0x000017bb-0x000017b8,1]}", -- 0x000017b8
    x"{code[0x000017bf-0x000017bc,1]}", -- 0x000017bc
    x"{code[0x000017c3-0x000017c0,1]}", -- 0x000017c0
    x"{code[0x000017c7-0x000017c4,1]}", -- 0x000017c4
    x"{code[0x000017cb-0x000017c8,1]}", -- 0x000017c8
    x"{code[0x000017cf-0x000017cc,1]}", -- 0x000017cc
    x"{code[0x000017d3-0x000017d0,1]}", -- 0x000017d0
    x"{code[0x000017d7-0x000017d4,1]}", -- 0x000017d4
    x"{code[0x000017db-0x000017d8,1]}", -- 0x000017d8
    x"{code[0x000017df-0x000017dc,1]}", -- 0x000017dc
    x"{code[0x000017e3-0x000017e0,1]}", -- 0x000017e0
    x"{code[0x000017e7-0x000017e4,1]}", -- 0x000017e4
    x"{code[0x000017eb-0x000017e8,1]}", -- 0x000017e8
    x"{code[0x000017ef-0x000017ec,1]}", -- 0x000017ec
    x"{code[0x000017f3-0x000017f0,1]}", -- 0x000017f0
    x"{code[0x000017f7-0x000017f4,1]}", -- 0x000017f4
    x"{code[0x000017fb-0x000017f8,1]}", -- 0x000017f8
    x"{code[0x000017ff-0x000017fc,1]}", -- 0x000017fc
    x"{code[0x00001803-0x00001800,1]}", -- 0x00001800
    x"{code[0x00001807-0x00001804,1]}", -- 0x00001804
    x"{code[0x0000180b-0x00001808,1]}", -- 0x00001808
    x"{code[0x0000180f-0x0000180c,1]}", -- 0x0000180c
    x"{code[0x00001813-0x00001810,1]}", -- 0x00001810
    x"{code[0x00001817-0x00001814,1]}", -- 0x00001814
    x"{code[0x0000181b-0x00001818,1]}", -- 0x00001818
    x"{code[0x0000181f-0x0000181c,1]}", -- 0x0000181c
    x"{code[0x00001823-0x00001820,1]}", -- 0x00001820
    x"{code[0x00001827-0x00001824,1]}", -- 0x00001824
    x"{code[0x0000182b-0x00001828,1]}", -- 0x00001828
    x"{code[0x0000182f-0x0000182c,1]}", -- 0x0000182c
    x"{code[0x00001833-0x00001830,1]}", -- 0x00001830
    x"{code[0x00001837-0x00001834,1]}", -- 0x00001834
    x"{code[0x0000183b-0x00001838,1]}", -- 0x00001838
    x"{code[0x0000183f-0x0000183c,1]}", -- 0x0000183c
    x"{code[0x00001843-0x00001840,1]}", -- 0x00001840
    x"{code[0x00001847-0x00001844,1]}", -- 0x00001844
    x"{code[0x0000184b-0x00001848,1]}", -- 0x00001848
    x"{code[0x0000184f-0x0000184c,1]}", -- 0x0000184c
    x"{code[0x00001853-0x00001850,1]}", -- 0x00001850
    x"{code[0x00001857-0x00001854,1]}", -- 0x00001854
    x"{code[0x0000185b-0x00001858,1]}", -- 0x00001858
    x"{code[0x0000185f-0x0000185c,1]}", -- 0x0000185c
    x"{code[0x00001863-0x00001860,1]}", -- 0x00001860
    x"{code[0x00001867-0x00001864,1]}", -- 0x00001864
    x"{code[0x0000186b-0x00001868,1]}", -- 0x00001868
    x"{code[0x0000186f-0x0000186c,1]}", -- 0x0000186c
    x"{code[0x00001873-0x00001870,1]}", -- 0x00001870
    x"{code[0x00001877-0x00001874,1]}", -- 0x00001874
    x"{code[0x0000187b-0x00001878,1]}", -- 0x00001878
    x"{code[0x0000187f-0x0000187c,1]}", -- 0x0000187c
    x"{code[0x00001883-0x00001880,1]}", -- 0x00001880
    x"{code[0x00001887-0x00001884,1]}", -- 0x00001884
    x"{code[0x0000188b-0x00001888,1]}", -- 0x00001888
    x"{code[0x0000188f-0x0000188c,1]}", -- 0x0000188c
    x"{code[0x00001893-0x00001890,1]}", -- 0x00001890
    x"{code[0x00001897-0x00001894,1]}", -- 0x00001894
    x"{code[0x0000189b-0x00001898,1]}", -- 0x00001898
    x"{code[0x0000189f-0x0000189c,1]}", -- 0x0000189c
    x"{code[0x000018a3-0x000018a0,1]}", -- 0x000018a0
    x"{code[0x000018a7-0x000018a4,1]}", -- 0x000018a4
    x"{code[0x000018ab-0x000018a8,1]}", -- 0x000018a8
    x"{code[0x000018af-0x000018ac,1]}", -- 0x000018ac
    x"{code[0x000018b3-0x000018b0,1]}", -- 0x000018b0
    x"{code[0x000018b7-0x000018b4,1]}", -- 0x000018b4
    x"{code[0x000018bb-0x000018b8,1]}", -- 0x000018b8
    x"{code[0x000018bf-0x000018bc,1]}", -- 0x000018bc
    x"{code[0x000018c3-0x000018c0,1]}", -- 0x000018c0
    x"{code[0x000018c7-0x000018c4,1]}", -- 0x000018c4
    x"{code[0x000018cb-0x000018c8,1]}", -- 0x000018c8
    x"{code[0x000018cf-0x000018cc,1]}", -- 0x000018cc
    x"{code[0x000018d3-0x000018d0,1]}", -- 0x000018d0
    x"{code[0x000018d7-0x000018d4,1]}", -- 0x000018d4
    x"{code[0x000018db-0x000018d8,1]}", -- 0x000018d8
    x"{code[0x000018df-0x000018dc,1]}", -- 0x000018dc
    x"{code[0x000018e3-0x000018e0,1]}", -- 0x000018e0
    x"{code[0x000018e7-0x000018e4,1]}", -- 0x000018e4
    x"{code[0x000018eb-0x000018e8,1]}", -- 0x000018e8
    x"{code[0x000018ef-0x000018ec,1]}", -- 0x000018ec
    x"{code[0x000018f3-0x000018f0,1]}", -- 0x000018f0
    x"{code[0x000018f7-0x000018f4,1]}", -- 0x000018f4
    x"{code[0x000018fb-0x000018f8,1]}", -- 0x000018f8
    x"{code[0x000018ff-0x000018fc,1]}", -- 0x000018fc
    x"{code[0x00001903-0x00001900,1]}", -- 0x00001900
    x"{code[0x00001907-0x00001904,1]}", -- 0x00001904
    x"{code[0x0000190b-0x00001908,1]}", -- 0x00001908
    x"{code[0x0000190f-0x0000190c,1]}", -- 0x0000190c
    x"{code[0x00001913-0x00001910,1]}", -- 0x00001910
    x"{code[0x00001917-0x00001914,1]}", -- 0x00001914
    x"{code[0x0000191b-0x00001918,1]}", -- 0x00001918
    x"{code[0x0000191f-0x0000191c,1]}", -- 0x0000191c
    x"{code[0x00001923-0x00001920,1]}", -- 0x00001920
    x"{code[0x00001927-0x00001924,1]}", -- 0x00001924
    x"{code[0x0000192b-0x00001928,1]}", -- 0x00001928
    x"{code[0x0000192f-0x0000192c,1]}", -- 0x0000192c
    x"{code[0x00001933-0x00001930,1]}", -- 0x00001930
    x"{code[0x00001937-0x00001934,1]}", -- 0x00001934
    x"{code[0x0000193b-0x00001938,1]}", -- 0x00001938
    x"{code[0x0000193f-0x0000193c,1]}", -- 0x0000193c
    x"{code[0x00001943-0x00001940,1]}", -- 0x00001940
    x"{code[0x00001947-0x00001944,1]}", -- 0x00001944
    x"{code[0x0000194b-0x00001948,1]}", -- 0x00001948
    x"{code[0x0000194f-0x0000194c,1]}", -- 0x0000194c
    x"{code[0x00001953-0x00001950,1]}", -- 0x00001950
    x"{code[0x00001957-0x00001954,1]}", -- 0x00001954
    x"{code[0x0000195b-0x00001958,1]}", -- 0x00001958
    x"{code[0x0000195f-0x0000195c,1]}", -- 0x0000195c
    x"{code[0x00001963-0x00001960,1]}", -- 0x00001960
    x"{code[0x00001967-0x00001964,1]}", -- 0x00001964
    x"{code[0x0000196b-0x00001968,1]}", -- 0x00001968
    x"{code[0x0000196f-0x0000196c,1]}", -- 0x0000196c
    x"{code[0x00001973-0x00001970,1]}", -- 0x00001970
    x"{code[0x00001977-0x00001974,1]}", -- 0x00001974
    x"{code[0x0000197b-0x00001978,1]}", -- 0x00001978
    x"{code[0x0000197f-0x0000197c,1]}", -- 0x0000197c
    x"{code[0x00001983-0x00001980,1]}", -- 0x00001980
    x"{code[0x00001987-0x00001984,1]}", -- 0x00001984
    x"{code[0x0000198b-0x00001988,1]}", -- 0x00001988
    x"{code[0x0000198f-0x0000198c,1]}", -- 0x0000198c
    x"{code[0x00001993-0x00001990,1]}", -- 0x00001990
    x"{code[0x00001997-0x00001994,1]}", -- 0x00001994
    x"{code[0x0000199b-0x00001998,1]}", -- 0x00001998
    x"{code[0x0000199f-0x0000199c,1]}", -- 0x0000199c
    x"{code[0x000019a3-0x000019a0,1]}", -- 0x000019a0
    x"{code[0x000019a7-0x000019a4,1]}", -- 0x000019a4
    x"{code[0x000019ab-0x000019a8,1]}", -- 0x000019a8
    x"{code[0x000019af-0x000019ac,1]}", -- 0x000019ac
    x"{code[0x000019b3-0x000019b0,1]}", -- 0x000019b0
    x"{code[0x000019b7-0x000019b4,1]}", -- 0x000019b4
    x"{code[0x000019bb-0x000019b8,1]}", -- 0x000019b8
    x"{code[0x000019bf-0x000019bc,1]}", -- 0x000019bc
    x"{code[0x000019c3-0x000019c0,1]}", -- 0x000019c0
    x"{code[0x000019c7-0x000019c4,1]}", -- 0x000019c4
    x"{code[0x000019cb-0x000019c8,1]}", -- 0x000019c8
    x"{code[0x000019cf-0x000019cc,1]}", -- 0x000019cc
    x"{code[0x000019d3-0x000019d0,1]}", -- 0x000019d0
    x"{code[0x000019d7-0x000019d4,1]}", -- 0x000019d4
    x"{code[0x000019db-0x000019d8,1]}", -- 0x000019d8
    x"{code[0x000019df-0x000019dc,1]}", -- 0x000019dc
    x"{code[0x000019e3-0x000019e0,1]}", -- 0x000019e0
    x"{code[0x000019e7-0x000019e4,1]}", -- 0x000019e4
    x"{code[0x000019eb-0x000019e8,1]}", -- 0x000019e8
    x"{code[0x000019ef-0x000019ec,1]}", -- 0x000019ec
    x"{code[0x000019f3-0x000019f0,1]}", -- 0x000019f0
    x"{code[0x000019f7-0x000019f4,1]}", -- 0x000019f4
    x"{code[0x000019fb-0x000019f8,1]}", -- 0x000019f8
    x"{code[0x000019ff-0x000019fc,1]}", -- 0x000019fc
    x"{code[0x00001a03-0x00001a00,1]}", -- 0x00001a00
    x"{code[0x00001a07-0x00001a04,1]}", -- 0x00001a04
    x"{code[0x00001a0b-0x00001a08,1]}", -- 0x00001a08
    x"{code[0x00001a0f-0x00001a0c,1]}", -- 0x00001a0c
    x"{code[0x00001a13-0x00001a10,1]}", -- 0x00001a10
    x"{code[0x00001a17-0x00001a14,1]}", -- 0x00001a14
    x"{code[0x00001a1b-0x00001a18,1]}", -- 0x00001a18
    x"{code[0x00001a1f-0x00001a1c,1]}", -- 0x00001a1c
    x"{code[0x00001a23-0x00001a20,1]}", -- 0x00001a20
    x"{code[0x00001a27-0x00001a24,1]}", -- 0x00001a24
    x"{code[0x00001a2b-0x00001a28,1]}", -- 0x00001a28
    x"{code[0x00001a2f-0x00001a2c,1]}", -- 0x00001a2c
    x"{code[0x00001a33-0x00001a30,1]}", -- 0x00001a30
    x"{code[0x00001a37-0x00001a34,1]}", -- 0x00001a34
    x"{code[0x00001a3b-0x00001a38,1]}", -- 0x00001a38
    x"{code[0x00001a3f-0x00001a3c,1]}", -- 0x00001a3c
    x"{code[0x00001a43-0x00001a40,1]}", -- 0x00001a40
    x"{code[0x00001a47-0x00001a44,1]}", -- 0x00001a44
    x"{code[0x00001a4b-0x00001a48,1]}", -- 0x00001a48
    x"{code[0x00001a4f-0x00001a4c,1]}", -- 0x00001a4c
    x"{code[0x00001a53-0x00001a50,1]}", -- 0x00001a50
    x"{code[0x00001a57-0x00001a54,1]}", -- 0x00001a54
    x"{code[0x00001a5b-0x00001a58,1]}", -- 0x00001a58
    x"{code[0x00001a5f-0x00001a5c,1]}", -- 0x00001a5c
    x"{code[0x00001a63-0x00001a60,1]}", -- 0x00001a60
    x"{code[0x00001a67-0x00001a64,1]}", -- 0x00001a64
    x"{code[0x00001a6b-0x00001a68,1]}", -- 0x00001a68
    x"{code[0x00001a6f-0x00001a6c,1]}", -- 0x00001a6c
    x"{code[0x00001a73-0x00001a70,1]}", -- 0x00001a70
    x"{code[0x00001a77-0x00001a74,1]}", -- 0x00001a74
    x"{code[0x00001a7b-0x00001a78,1]}", -- 0x00001a78
    x"{code[0x00001a7f-0x00001a7c,1]}", -- 0x00001a7c
    x"{code[0x00001a83-0x00001a80,1]}", -- 0x00001a80
    x"{code[0x00001a87-0x00001a84,1]}", -- 0x00001a84
    x"{code[0x00001a8b-0x00001a88,1]}", -- 0x00001a88
    x"{code[0x00001a8f-0x00001a8c,1]}", -- 0x00001a8c
    x"{code[0x00001a93-0x00001a90,1]}", -- 0x00001a90
    x"{code[0x00001a97-0x00001a94,1]}", -- 0x00001a94
    x"{code[0x00001a9b-0x00001a98,1]}", -- 0x00001a98
    x"{code[0x00001a9f-0x00001a9c,1]}", -- 0x00001a9c
    x"{code[0x00001aa3-0x00001aa0,1]}", -- 0x00001aa0
    x"{code[0x00001aa7-0x00001aa4,1]}", -- 0x00001aa4
    x"{code[0x00001aab-0x00001aa8,1]}", -- 0x00001aa8
    x"{code[0x00001aaf-0x00001aac,1]}", -- 0x00001aac
    x"{code[0x00001ab3-0x00001ab0,1]}", -- 0x00001ab0
    x"{code[0x00001ab7-0x00001ab4,1]}", -- 0x00001ab4
    x"{code[0x00001abb-0x00001ab8,1]}", -- 0x00001ab8
    x"{code[0x00001abf-0x00001abc,1]}", -- 0x00001abc
    x"{code[0x00001ac3-0x00001ac0,1]}", -- 0x00001ac0
    x"{code[0x00001ac7-0x00001ac4,1]}", -- 0x00001ac4
    x"{code[0x00001acb-0x00001ac8,1]}", -- 0x00001ac8
    x"{code[0x00001acf-0x00001acc,1]}", -- 0x00001acc
    x"{code[0x00001ad3-0x00001ad0,1]}", -- 0x00001ad0
    x"{code[0x00001ad7-0x00001ad4,1]}", -- 0x00001ad4
    x"{code[0x00001adb-0x00001ad8,1]}", -- 0x00001ad8
    x"{code[0x00001adf-0x00001adc,1]}", -- 0x00001adc
    x"{code[0x00001ae3-0x00001ae0,1]}", -- 0x00001ae0
    x"{code[0x00001ae7-0x00001ae4,1]}", -- 0x00001ae4
    x"{code[0x00001aeb-0x00001ae8,1]}", -- 0x00001ae8
    x"{code[0x00001aef-0x00001aec,1]}", -- 0x00001aec
    x"{code[0x00001af3-0x00001af0,1]}", -- 0x00001af0
    x"{code[0x00001af7-0x00001af4,1]}", -- 0x00001af4
    x"{code[0x00001afb-0x00001af8,1]}", -- 0x00001af8
    x"{code[0x00001aff-0x00001afc,1]}", -- 0x00001afc
    x"{code[0x00001b03-0x00001b00,1]}", -- 0x00001b00
    x"{code[0x00001b07-0x00001b04,1]}", -- 0x00001b04
    x"{code[0x00001b0b-0x00001b08,1]}", -- 0x00001b08
    x"{code[0x00001b0f-0x00001b0c,1]}", -- 0x00001b0c
    x"{code[0x00001b13-0x00001b10,1]}", -- 0x00001b10
    x"{code[0x00001b17-0x00001b14,1]}", -- 0x00001b14
    x"{code[0x00001b1b-0x00001b18,1]}", -- 0x00001b18
    x"{code[0x00001b1f-0x00001b1c,1]}", -- 0x00001b1c
    x"{code[0x00001b23-0x00001b20,1]}", -- 0x00001b20
    x"{code[0x00001b27-0x00001b24,1]}", -- 0x00001b24
    x"{code[0x00001b2b-0x00001b28,1]}", -- 0x00001b28
    x"{code[0x00001b2f-0x00001b2c,1]}", -- 0x00001b2c
    x"{code[0x00001b33-0x00001b30,1]}", -- 0x00001b30
    x"{code[0x00001b37-0x00001b34,1]}", -- 0x00001b34
    x"{code[0x00001b3b-0x00001b38,1]}", -- 0x00001b38
    x"{code[0x00001b3f-0x00001b3c,1]}", -- 0x00001b3c
    x"{code[0x00001b43-0x00001b40,1]}", -- 0x00001b40
    x"{code[0x00001b47-0x00001b44,1]}", -- 0x00001b44
    x"{code[0x00001b4b-0x00001b48,1]}", -- 0x00001b48
    x"{code[0x00001b4f-0x00001b4c,1]}", -- 0x00001b4c
    x"{code[0x00001b53-0x00001b50,1]}", -- 0x00001b50
    x"{code[0x00001b57-0x00001b54,1]}", -- 0x00001b54
    x"{code[0x00001b5b-0x00001b58,1]}", -- 0x00001b58
    x"{code[0x00001b5f-0x00001b5c,1]}", -- 0x00001b5c
    x"{code[0x00001b63-0x00001b60,1]}", -- 0x00001b60
    x"{code[0x00001b67-0x00001b64,1]}", -- 0x00001b64
    x"{code[0x00001b6b-0x00001b68,1]}", -- 0x00001b68
    x"{code[0x00001b6f-0x00001b6c,1]}", -- 0x00001b6c
    x"{code[0x00001b73-0x00001b70,1]}", -- 0x00001b70
    x"{code[0x00001b77-0x00001b74,1]}", -- 0x00001b74
    x"{code[0x00001b7b-0x00001b78,1]}", -- 0x00001b78
    x"{code[0x00001b7f-0x00001b7c,1]}", -- 0x00001b7c
    x"{code[0x00001b83-0x00001b80,1]}", -- 0x00001b80
    x"{code[0x00001b87-0x00001b84,1]}", -- 0x00001b84
    x"{code[0x00001b8b-0x00001b88,1]}", -- 0x00001b88
    x"{code[0x00001b8f-0x00001b8c,1]}", -- 0x00001b8c
    x"{code[0x00001b93-0x00001b90,1]}", -- 0x00001b90
    x"{code[0x00001b97-0x00001b94,1]}", -- 0x00001b94
    x"{code[0x00001b9b-0x00001b98,1]}", -- 0x00001b98
    x"{code[0x00001b9f-0x00001b9c,1]}", -- 0x00001b9c
    x"{code[0x00001ba3-0x00001ba0,1]}", -- 0x00001ba0
    x"{code[0x00001ba7-0x00001ba4,1]}", -- 0x00001ba4
    x"{code[0x00001bab-0x00001ba8,1]}", -- 0x00001ba8
    x"{code[0x00001baf-0x00001bac,1]}", -- 0x00001bac
    x"{code[0x00001bb3-0x00001bb0,1]}", -- 0x00001bb0
    x"{code[0x00001bb7-0x00001bb4,1]}", -- 0x00001bb4
    x"{code[0x00001bbb-0x00001bb8,1]}", -- 0x00001bb8
    x"{code[0x00001bbf-0x00001bbc,1]}", -- 0x00001bbc
    x"{code[0x00001bc3-0x00001bc0,1]}", -- 0x00001bc0
    x"{code[0x00001bc7-0x00001bc4,1]}", -- 0x00001bc4
    x"{code[0x00001bcb-0x00001bc8,1]}", -- 0x00001bc8
    x"{code[0x00001bcf-0x00001bcc,1]}", -- 0x00001bcc
    x"{code[0x00001bd3-0x00001bd0,1]}", -- 0x00001bd0
    x"{code[0x00001bd7-0x00001bd4,1]}", -- 0x00001bd4
    x"{code[0x00001bdb-0x00001bd8,1]}", -- 0x00001bd8
    x"{code[0x00001bdf-0x00001bdc,1]}", -- 0x00001bdc
    x"{code[0x00001be3-0x00001be0,1]}", -- 0x00001be0
    x"{code[0x00001be7-0x00001be4,1]}", -- 0x00001be4
    x"{code[0x00001beb-0x00001be8,1]}", -- 0x00001be8
    x"{code[0x00001bef-0x00001bec,1]}", -- 0x00001bec
    x"{code[0x00001bf3-0x00001bf0,1]}", -- 0x00001bf0
    x"{code[0x00001bf7-0x00001bf4,1]}", -- 0x00001bf4
    x"{code[0x00001bfb-0x00001bf8,1]}", -- 0x00001bf8
    x"{code[0x00001bff-0x00001bfc,1]}", -- 0x00001bfc
    x"{code[0x00001c03-0x00001c00,1]}", -- 0x00001c00
    x"{code[0x00001c07-0x00001c04,1]}", -- 0x00001c04
    x"{code[0x00001c0b-0x00001c08,1]}", -- 0x00001c08
    x"{code[0x00001c0f-0x00001c0c,1]}", -- 0x00001c0c
    x"{code[0x00001c13-0x00001c10,1]}", -- 0x00001c10
    x"{code[0x00001c17-0x00001c14,1]}", -- 0x00001c14
    x"{code[0x00001c1b-0x00001c18,1]}", -- 0x00001c18
    x"{code[0x00001c1f-0x00001c1c,1]}", -- 0x00001c1c
    x"{code[0x00001c23-0x00001c20,1]}", -- 0x00001c20
    x"{code[0x00001c27-0x00001c24,1]}", -- 0x00001c24
    x"{code[0x00001c2b-0x00001c28,1]}", -- 0x00001c28
    x"{code[0x00001c2f-0x00001c2c,1]}", -- 0x00001c2c
    x"{code[0x00001c33-0x00001c30,1]}", -- 0x00001c30
    x"{code[0x00001c37-0x00001c34,1]}", -- 0x00001c34
    x"{code[0x00001c3b-0x00001c38,1]}", -- 0x00001c38
    x"{code[0x00001c3f-0x00001c3c,1]}", -- 0x00001c3c
    x"{code[0x00001c43-0x00001c40,1]}", -- 0x00001c40
    x"{code[0x00001c47-0x00001c44,1]}", -- 0x00001c44
    x"{code[0x00001c4b-0x00001c48,1]}", -- 0x00001c48
    x"{code[0x00001c4f-0x00001c4c,1]}", -- 0x00001c4c
    x"{code[0x00001c53-0x00001c50,1]}", -- 0x00001c50
    x"{code[0x00001c57-0x00001c54,1]}", -- 0x00001c54
    x"{code[0x00001c5b-0x00001c58,1]}", -- 0x00001c58
    x"{code[0x00001c5f-0x00001c5c,1]}", -- 0x00001c5c
    x"{code[0x00001c63-0x00001c60,1]}", -- 0x00001c60
    x"{code[0x00001c67-0x00001c64,1]}", -- 0x00001c64
    x"{code[0x00001c6b-0x00001c68,1]}", -- 0x00001c68
    x"{code[0x00001c6f-0x00001c6c,1]}", -- 0x00001c6c
    x"{code[0x00001c73-0x00001c70,1]}", -- 0x00001c70
    x"{code[0x00001c77-0x00001c74,1]}", -- 0x00001c74
    x"{code[0x00001c7b-0x00001c78,1]}", -- 0x00001c78
    x"{code[0x00001c7f-0x00001c7c,1]}", -- 0x00001c7c
    x"{code[0x00001c83-0x00001c80,1]}", -- 0x00001c80
    x"{code[0x00001c87-0x00001c84,1]}", -- 0x00001c84
    x"{code[0x00001c8b-0x00001c88,1]}", -- 0x00001c88
    x"{code[0x00001c8f-0x00001c8c,1]}", -- 0x00001c8c
    x"{code[0x00001c93-0x00001c90,1]}", -- 0x00001c90
    x"{code[0x00001c97-0x00001c94,1]}", -- 0x00001c94
    x"{code[0x00001c9b-0x00001c98,1]}", -- 0x00001c98
    x"{code[0x00001c9f-0x00001c9c,1]}", -- 0x00001c9c
    x"{code[0x00001ca3-0x00001ca0,1]}", -- 0x00001ca0
    x"{code[0x00001ca7-0x00001ca4,1]}", -- 0x00001ca4
    x"{code[0x00001cab-0x00001ca8,1]}", -- 0x00001ca8
    x"{code[0x00001caf-0x00001cac,1]}", -- 0x00001cac
    x"{code[0x00001cb3-0x00001cb0,1]}", -- 0x00001cb0
    x"{code[0x00001cb7-0x00001cb4,1]}", -- 0x00001cb4
    x"{code[0x00001cbb-0x00001cb8,1]}", -- 0x00001cb8
    x"{code[0x00001cbf-0x00001cbc,1]}", -- 0x00001cbc
    x"{code[0x00001cc3-0x00001cc0,1]}", -- 0x00001cc0
    x"{code[0x00001cc7-0x00001cc4,1]}", -- 0x00001cc4
    x"{code[0x00001ccb-0x00001cc8,1]}", -- 0x00001cc8
    x"{code[0x00001ccf-0x00001ccc,1]}", -- 0x00001ccc
    x"{code[0x00001cd3-0x00001cd0,1]}", -- 0x00001cd0
    x"{code[0x00001cd7-0x00001cd4,1]}", -- 0x00001cd4
    x"{code[0x00001cdb-0x00001cd8,1]}", -- 0x00001cd8
    x"{code[0x00001cdf-0x00001cdc,1]}", -- 0x00001cdc
    x"{code[0x00001ce3-0x00001ce0,1]}", -- 0x00001ce0
    x"{code[0x00001ce7-0x00001ce4,1]}", -- 0x00001ce4
    x"{code[0x00001ceb-0x00001ce8,1]}", -- 0x00001ce8
    x"{code[0x00001cef-0x00001cec,1]}", -- 0x00001cec
    x"{code[0x00001cf3-0x00001cf0,1]}", -- 0x00001cf0
    x"{code[0x00001cf7-0x00001cf4,1]}", -- 0x00001cf4
    x"{code[0x00001cfb-0x00001cf8,1]}", -- 0x00001cf8
    x"{code[0x00001cff-0x00001cfc,1]}", -- 0x00001cfc
    x"{code[0x00001d03-0x00001d00,1]}", -- 0x00001d00
    x"{code[0x00001d07-0x00001d04,1]}", -- 0x00001d04
    x"{code[0x00001d0b-0x00001d08,1]}", -- 0x00001d08
    x"{code[0x00001d0f-0x00001d0c,1]}", -- 0x00001d0c
    x"{code[0x00001d13-0x00001d10,1]}", -- 0x00001d10
    x"{code[0x00001d17-0x00001d14,1]}", -- 0x00001d14
    x"{code[0x00001d1b-0x00001d18,1]}", -- 0x00001d18
    x"{code[0x00001d1f-0x00001d1c,1]}", -- 0x00001d1c
    x"{code[0x00001d23-0x00001d20,1]}", -- 0x00001d20
    x"{code[0x00001d27-0x00001d24,1]}", -- 0x00001d24
    x"{code[0x00001d2b-0x00001d28,1]}", -- 0x00001d28
    x"{code[0x00001d2f-0x00001d2c,1]}", -- 0x00001d2c
    x"{code[0x00001d33-0x00001d30,1]}", -- 0x00001d30
    x"{code[0x00001d37-0x00001d34,1]}", -- 0x00001d34
    x"{code[0x00001d3b-0x00001d38,1]}", -- 0x00001d38
    x"{code[0x00001d3f-0x00001d3c,1]}", -- 0x00001d3c
    x"{code[0x00001d43-0x00001d40,1]}", -- 0x00001d40
    x"{code[0x00001d47-0x00001d44,1]}", -- 0x00001d44
    x"{code[0x00001d4b-0x00001d48,1]}", -- 0x00001d48
    x"{code[0x00001d4f-0x00001d4c,1]}", -- 0x00001d4c
    x"{code[0x00001d53-0x00001d50,1]}", -- 0x00001d50
    x"{code[0x00001d57-0x00001d54,1]}", -- 0x00001d54
    x"{code[0x00001d5b-0x00001d58,1]}", -- 0x00001d58
    x"{code[0x00001d5f-0x00001d5c,1]}", -- 0x00001d5c
    x"{code[0x00001d63-0x00001d60,1]}", -- 0x00001d60
    x"{code[0x00001d67-0x00001d64,1]}", -- 0x00001d64
    x"{code[0x00001d6b-0x00001d68,1]}", -- 0x00001d68
    x"{code[0x00001d6f-0x00001d6c,1]}", -- 0x00001d6c
    x"{code[0x00001d73-0x00001d70,1]}", -- 0x00001d70
    x"{code[0x00001d77-0x00001d74,1]}", -- 0x00001d74
    x"{code[0x00001d7b-0x00001d78,1]}", -- 0x00001d78
    x"{code[0x00001d7f-0x00001d7c,1]}", -- 0x00001d7c
    x"{code[0x00001d83-0x00001d80,1]}", -- 0x00001d80
    x"{code[0x00001d87-0x00001d84,1]}", -- 0x00001d84
    x"{code[0x00001d8b-0x00001d88,1]}", -- 0x00001d88
    x"{code[0x00001d8f-0x00001d8c,1]}", -- 0x00001d8c
    x"{code[0x00001d93-0x00001d90,1]}", -- 0x00001d90
    x"{code[0x00001d97-0x00001d94,1]}", -- 0x00001d94
    x"{code[0x00001d9b-0x00001d98,1]}", -- 0x00001d98
    x"{code[0x00001d9f-0x00001d9c,1]}", -- 0x00001d9c
    x"{code[0x00001da3-0x00001da0,1]}", -- 0x00001da0
    x"{code[0x00001da7-0x00001da4,1]}", -- 0x00001da4
    x"{code[0x00001dab-0x00001da8,1]}", -- 0x00001da8
    x"{code[0x00001daf-0x00001dac,1]}", -- 0x00001dac
    x"{code[0x00001db3-0x00001db0,1]}", -- 0x00001db0
    x"{code[0x00001db7-0x00001db4,1]}", -- 0x00001db4
    x"{code[0x00001dbb-0x00001db8,1]}", -- 0x00001db8
    x"{code[0x00001dbf-0x00001dbc,1]}", -- 0x00001dbc
    x"{code[0x00001dc3-0x00001dc0,1]}", -- 0x00001dc0
    x"{code[0x00001dc7-0x00001dc4,1]}", -- 0x00001dc4
    x"{code[0x00001dcb-0x00001dc8,1]}", -- 0x00001dc8
    x"{code[0x00001dcf-0x00001dcc,1]}", -- 0x00001dcc
    x"{code[0x00001dd3-0x00001dd0,1]}", -- 0x00001dd0
    x"{code[0x00001dd7-0x00001dd4,1]}", -- 0x00001dd4
    x"{code[0x00001ddb-0x00001dd8,1]}", -- 0x00001dd8
    x"{code[0x00001ddf-0x00001ddc,1]}", -- 0x00001ddc
    x"{code[0x00001de3-0x00001de0,1]}", -- 0x00001de0
    x"{code[0x00001de7-0x00001de4,1]}", -- 0x00001de4
    x"{code[0x00001deb-0x00001de8,1]}", -- 0x00001de8
    x"{code[0x00001def-0x00001dec,1]}", -- 0x00001dec
    x"{code[0x00001df3-0x00001df0,1]}", -- 0x00001df0
    x"{code[0x00001df7-0x00001df4,1]}", -- 0x00001df4
    x"{code[0x00001dfb-0x00001df8,1]}", -- 0x00001df8
    x"{code[0x00001dff-0x00001dfc,1]}", -- 0x00001dfc
    x"{code[0x00001e03-0x00001e00,1]}", -- 0x00001e00
    x"{code[0x00001e07-0x00001e04,1]}", -- 0x00001e04
    x"{code[0x00001e0b-0x00001e08,1]}", -- 0x00001e08
    x"{code[0x00001e0f-0x00001e0c,1]}", -- 0x00001e0c
    x"{code[0x00001e13-0x00001e10,1]}", -- 0x00001e10
    x"{code[0x00001e17-0x00001e14,1]}", -- 0x00001e14
    x"{code[0x00001e1b-0x00001e18,1]}", -- 0x00001e18
    x"{code[0x00001e1f-0x00001e1c,1]}", -- 0x00001e1c
    x"{code[0x00001e23-0x00001e20,1]}", -- 0x00001e20
    x"{code[0x00001e27-0x00001e24,1]}", -- 0x00001e24
    x"{code[0x00001e2b-0x00001e28,1]}", -- 0x00001e28
    x"{code[0x00001e2f-0x00001e2c,1]}", -- 0x00001e2c
    x"{code[0x00001e33-0x00001e30,1]}", -- 0x00001e30
    x"{code[0x00001e37-0x00001e34,1]}", -- 0x00001e34
    x"{code[0x00001e3b-0x00001e38,1]}", -- 0x00001e38
    x"{code[0x00001e3f-0x00001e3c,1]}", -- 0x00001e3c
    x"{code[0x00001e43-0x00001e40,1]}", -- 0x00001e40
    x"{code[0x00001e47-0x00001e44,1]}", -- 0x00001e44
    x"{code[0x00001e4b-0x00001e48,1]}", -- 0x00001e48
    x"{code[0x00001e4f-0x00001e4c,1]}", -- 0x00001e4c
    x"{code[0x00001e53-0x00001e50,1]}", -- 0x00001e50
    x"{code[0x00001e57-0x00001e54,1]}", -- 0x00001e54
    x"{code[0x00001e5b-0x00001e58,1]}", -- 0x00001e58
    x"{code[0x00001e5f-0x00001e5c,1]}", -- 0x00001e5c
    x"{code[0x00001e63-0x00001e60,1]}", -- 0x00001e60
    x"{code[0x00001e67-0x00001e64,1]}", -- 0x00001e64
    x"{code[0x00001e6b-0x00001e68,1]}", -- 0x00001e68
    x"{code[0x00001e6f-0x00001e6c,1]}", -- 0x00001e6c
    x"{code[0x00001e73-0x00001e70,1]}", -- 0x00001e70
    x"{code[0x00001e77-0x00001e74,1]}", -- 0x00001e74
    x"{code[0x00001e7b-0x00001e78,1]}", -- 0x00001e78
    x"{code[0x00001e7f-0x00001e7c,1]}", -- 0x00001e7c
    x"{code[0x00001e83-0x00001e80,1]}", -- 0x00001e80
    x"{code[0x00001e87-0x00001e84,1]}", -- 0x00001e84
    x"{code[0x00001e8b-0x00001e88,1]}", -- 0x00001e88
    x"{code[0x00001e8f-0x00001e8c,1]}", -- 0x00001e8c
    x"{code[0x00001e93-0x00001e90,1]}", -- 0x00001e90
    x"{code[0x00001e97-0x00001e94,1]}", -- 0x00001e94
    x"{code[0x00001e9b-0x00001e98,1]}", -- 0x00001e98
    x"{code[0x00001e9f-0x00001e9c,1]}", -- 0x00001e9c
    x"{code[0x00001ea3-0x00001ea0,1]}", -- 0x00001ea0
    x"{code[0x00001ea7-0x00001ea4,1]}", -- 0x00001ea4
    x"{code[0x00001eab-0x00001ea8,1]}", -- 0x00001ea8
    x"{code[0x00001eaf-0x00001eac,1]}", -- 0x00001eac
    x"{code[0x00001eb3-0x00001eb0,1]}", -- 0x00001eb0
    x"{code[0x00001eb7-0x00001eb4,1]}", -- 0x00001eb4
    x"{code[0x00001ebb-0x00001eb8,1]}", -- 0x00001eb8
    x"{code[0x00001ebf-0x00001ebc,1]}", -- 0x00001ebc
    x"{code[0x00001ec3-0x00001ec0,1]}", -- 0x00001ec0
    x"{code[0x00001ec7-0x00001ec4,1]}", -- 0x00001ec4
    x"{code[0x00001ecb-0x00001ec8,1]}", -- 0x00001ec8
    x"{code[0x00001ecf-0x00001ecc,1]}", -- 0x00001ecc
    x"{code[0x00001ed3-0x00001ed0,1]}", -- 0x00001ed0
    x"{code[0x00001ed7-0x00001ed4,1]}", -- 0x00001ed4
    x"{code[0x00001edb-0x00001ed8,1]}", -- 0x00001ed8
    x"{code[0x00001edf-0x00001edc,1]}", -- 0x00001edc
    x"{code[0x00001ee3-0x00001ee0,1]}", -- 0x00001ee0
    x"{code[0x00001ee7-0x00001ee4,1]}", -- 0x00001ee4
    x"{code[0x00001eeb-0x00001ee8,1]}", -- 0x00001ee8
    x"{code[0x00001eef-0x00001eec,1]}", -- 0x00001eec
    x"{code[0x00001ef3-0x00001ef0,1]}", -- 0x00001ef0
    x"{code[0x00001ef7-0x00001ef4,1]}", -- 0x00001ef4
    x"{code[0x00001efb-0x00001ef8,1]}", -- 0x00001ef8
    x"{code[0x00001eff-0x00001efc,1]}", -- 0x00001efc
    x"{code[0x00001f03-0x00001f00,1]}", -- 0x00001f00
    x"{code[0x00001f07-0x00001f04,1]}", -- 0x00001f04
    x"{code[0x00001f0b-0x00001f08,1]}", -- 0x00001f08
    x"{code[0x00001f0f-0x00001f0c,1]}", -- 0x00001f0c
    x"{code[0x00001f13-0x00001f10,1]}", -- 0x00001f10
    x"{code[0x00001f17-0x00001f14,1]}", -- 0x00001f14
    x"{code[0x00001f1b-0x00001f18,1]}", -- 0x00001f18
    x"{code[0x00001f1f-0x00001f1c,1]}", -- 0x00001f1c
    x"{code[0x00001f23-0x00001f20,1]}", -- 0x00001f20
    x"{code[0x00001f27-0x00001f24,1]}", -- 0x00001f24
    x"{code[0x00001f2b-0x00001f28,1]}", -- 0x00001f28
    x"{code[0x00001f2f-0x00001f2c,1]}", -- 0x00001f2c
    x"{code[0x00001f33-0x00001f30,1]}", -- 0x00001f30
    x"{code[0x00001f37-0x00001f34,1]}", -- 0x00001f34
    x"{code[0x00001f3b-0x00001f38,1]}", -- 0x00001f38
    x"{code[0x00001f3f-0x00001f3c,1]}", -- 0x00001f3c
    x"{code[0x00001f43-0x00001f40,1]}", -- 0x00001f40
    x"{code[0x00001f47-0x00001f44,1]}", -- 0x00001f44
    x"{code[0x00001f4b-0x00001f48,1]}", -- 0x00001f48
    x"{code[0x00001f4f-0x00001f4c,1]}", -- 0x00001f4c
    x"{code[0x00001f53-0x00001f50,1]}", -- 0x00001f50
    x"{code[0x00001f57-0x00001f54,1]}", -- 0x00001f54
    x"{code[0x00001f5b-0x00001f58,1]}", -- 0x00001f58
    x"{code[0x00001f5f-0x00001f5c,1]}", -- 0x00001f5c
    x"{code[0x00001f63-0x00001f60,1]}", -- 0x00001f60
    x"{code[0x00001f67-0x00001f64,1]}", -- 0x00001f64
    x"{code[0x00001f6b-0x00001f68,1]}", -- 0x00001f68
    x"{code[0x00001f6f-0x00001f6c,1]}", -- 0x00001f6c
    x"{code[0x00001f73-0x00001f70,1]}", -- 0x00001f70
    x"{code[0x00001f77-0x00001f74,1]}", -- 0x00001f74
    x"{code[0x00001f7b-0x00001f78,1]}", -- 0x00001f78
    x"{code[0x00001f7f-0x00001f7c,1]}", -- 0x00001f7c
    x"{code[0x00001f83-0x00001f80,1]}", -- 0x00001f80
    x"{code[0x00001f87-0x00001f84,1]}", -- 0x00001f84
    x"{code[0x00001f8b-0x00001f88,1]}", -- 0x00001f88
    x"{code[0x00001f8f-0x00001f8c,1]}", -- 0x00001f8c
    x"{code[0x00001f93-0x00001f90,1]}", -- 0x00001f90
    x"{code[0x00001f97-0x00001f94,1]}", -- 0x00001f94
    x"{code[0x00001f9b-0x00001f98,1]}", -- 0x00001f98
    x"{code[0x00001f9f-0x00001f9c,1]}", -- 0x00001f9c
    x"{code[0x00001fa3-0x00001fa0,1]}", -- 0x00001fa0
    x"{code[0x00001fa7-0x00001fa4,1]}", -- 0x00001fa4
    x"{code[0x00001fab-0x00001fa8,1]}", -- 0x00001fa8
    x"{code[0x00001faf-0x00001fac,1]}", -- 0x00001fac
    x"{code[0x00001fb3-0x00001fb0,1]}", -- 0x00001fb0
    x"{code[0x00001fb7-0x00001fb4,1]}", -- 0x00001fb4
    x"{code[0x00001fbb-0x00001fb8,1]}", -- 0x00001fb8
    x"{code[0x00001fbf-0x00001fbc,1]}", -- 0x00001fbc
    x"{code[0x00001fc3-0x00001fc0,1]}", -- 0x00001fc0
    x"{code[0x00001fc7-0x00001fc4,1]}", -- 0x00001fc4
    x"{code[0x00001fcb-0x00001fc8,1]}", -- 0x00001fc8
    x"{code[0x00001fcf-0x00001fcc,1]}", -- 0x00001fcc
    x"{code[0x00001fd3-0x00001fd0,1]}", -- 0x00001fd0
    x"{code[0x00001fd7-0x00001fd4,1]}", -- 0x00001fd4
    x"{code[0x00001fdb-0x00001fd8,1]}", -- 0x00001fd8
    x"{code[0x00001fdf-0x00001fdc,1]}", -- 0x00001fdc
    x"{code[0x00001fe3-0x00001fe0,1]}", -- 0x00001fe0
    x"{code[0x00001fe7-0x00001fe4,1]}", -- 0x00001fe4
    x"{code[0x00001feb-0x00001fe8,1]}", -- 0x00001fe8
    x"{code[0x00001fef-0x00001fec,1]}", -- 0x00001fec
    x"{code[0x00001ff3-0x00001ff0,1]}", -- 0x00001ff0
    x"{code[0x00001ff7-0x00001ff4,1]}", -- 0x00001ff4
    x"{code[0x00001ffb-0x00001ff8,1]}", -- 0x00001ff8
    x"{code[0x00001fff-0x00001ffc,1]}", -- 0x00001ffc
    x"{code[0x00002003-0x00002000,1]}", -- 0x00002000
    x"{code[0x00002007-0x00002004,1]}", -- 0x00002004
    x"{code[0x0000200b-0x00002008,1]}", -- 0x00002008
    x"{code[0x0000200f-0x0000200c,1]}", -- 0x0000200c
    x"{code[0x00002013-0x00002010,1]}", -- 0x00002010
    x"{code[0x00002017-0x00002014,1]}", -- 0x00002014
    x"{code[0x0000201b-0x00002018,1]}", -- 0x00002018
    x"{code[0x0000201f-0x0000201c,1]}", -- 0x0000201c
    x"{code[0x00002023-0x00002020,1]}", -- 0x00002020
    x"{code[0x00002027-0x00002024,1]}", -- 0x00002024
    x"{code[0x0000202b-0x00002028,1]}", -- 0x00002028
    x"{code[0x0000202f-0x0000202c,1]}", -- 0x0000202c
    x"{code[0x00002033-0x00002030,1]}", -- 0x00002030
    x"{code[0x00002037-0x00002034,1]}", -- 0x00002034
    x"{code[0x0000203b-0x00002038,1]}", -- 0x00002038
    x"{code[0x0000203f-0x0000203c,1]}", -- 0x0000203c
    x"{code[0x00002043-0x00002040,1]}", -- 0x00002040
    x"{code[0x00002047-0x00002044,1]}", -- 0x00002044
    x"{code[0x0000204b-0x00002048,1]}", -- 0x00002048
    x"{code[0x0000204f-0x0000204c,1]}", -- 0x0000204c
    x"{code[0x00002053-0x00002050,1]}", -- 0x00002050
    x"{code[0x00002057-0x00002054,1]}", -- 0x00002054
    x"{code[0x0000205b-0x00002058,1]}", -- 0x00002058
    x"{code[0x0000205f-0x0000205c,1]}", -- 0x0000205c
    x"{code[0x00002063-0x00002060,1]}", -- 0x00002060
    x"{code[0x00002067-0x00002064,1]}", -- 0x00002064
    x"{code[0x0000206b-0x00002068,1]}", -- 0x00002068
    x"{code[0x0000206f-0x0000206c,1]}", -- 0x0000206c
    x"{code[0x00002073-0x00002070,1]}", -- 0x00002070
    x"{code[0x00002077-0x00002074,1]}", -- 0x00002074
    x"{code[0x0000207b-0x00002078,1]}", -- 0x00002078
    x"{code[0x0000207f-0x0000207c,1]}", -- 0x0000207c
    x"{code[0x00002083-0x00002080,1]}", -- 0x00002080
    x"{code[0x00002087-0x00002084,1]}", -- 0x00002084
    x"{code[0x0000208b-0x00002088,1]}", -- 0x00002088
    x"{code[0x0000208f-0x0000208c,1]}", -- 0x0000208c
    x"{code[0x00002093-0x00002090,1]}", -- 0x00002090
    x"{code[0x00002097-0x00002094,1]}", -- 0x00002094
    x"{code[0x0000209b-0x00002098,1]}", -- 0x00002098
    x"{code[0x0000209f-0x0000209c,1]}", -- 0x0000209c
    x"{code[0x000020a3-0x000020a0,1]}", -- 0x000020a0
    x"{code[0x000020a7-0x000020a4,1]}", -- 0x000020a4
    x"{code[0x000020ab-0x000020a8,1]}", -- 0x000020a8
    x"{code[0x000020af-0x000020ac,1]}", -- 0x000020ac
    x"{code[0x000020b3-0x000020b0,1]}", -- 0x000020b0
    x"{code[0x000020b7-0x000020b4,1]}", -- 0x000020b4
    x"{code[0x000020bb-0x000020b8,1]}", -- 0x000020b8
    x"{code[0x000020bf-0x000020bc,1]}", -- 0x000020bc
    x"{code[0x000020c3-0x000020c0,1]}", -- 0x000020c0
    x"{code[0x000020c7-0x000020c4,1]}", -- 0x000020c4
    x"{code[0x000020cb-0x000020c8,1]}", -- 0x000020c8
    x"{code[0x000020cf-0x000020cc,1]}", -- 0x000020cc
    x"{code[0x000020d3-0x000020d0,1]}", -- 0x000020d0
    x"{code[0x000020d7-0x000020d4,1]}", -- 0x000020d4
    x"{code[0x000020db-0x000020d8,1]}", -- 0x000020d8
    x"{code[0x000020df-0x000020dc,1]}", -- 0x000020dc
    x"{code[0x000020e3-0x000020e0,1]}", -- 0x000020e0
    x"{code[0x000020e7-0x000020e4,1]}", -- 0x000020e4
    x"{code[0x000020eb-0x000020e8,1]}", -- 0x000020e8
    x"{code[0x000020ef-0x000020ec,1]}", -- 0x000020ec
    x"{code[0x000020f3-0x000020f0,1]}", -- 0x000020f0
    x"{code[0x000020f7-0x000020f4,1]}", -- 0x000020f4
    x"{code[0x000020fb-0x000020f8,1]}", -- 0x000020f8
    x"{code[0x000020ff-0x000020fc,1]}", -- 0x000020fc
    x"{code[0x00002103-0x00002100,1]}", -- 0x00002100
    x"{code[0x00002107-0x00002104,1]}", -- 0x00002104
    x"{code[0x0000210b-0x00002108,1]}", -- 0x00002108
    x"{code[0x0000210f-0x0000210c,1]}", -- 0x0000210c
    x"{code[0x00002113-0x00002110,1]}", -- 0x00002110
    x"{code[0x00002117-0x00002114,1]}", -- 0x00002114
    x"{code[0x0000211b-0x00002118,1]}", -- 0x00002118
    x"{code[0x0000211f-0x0000211c,1]}", -- 0x0000211c
    x"{code[0x00002123-0x00002120,1]}", -- 0x00002120
    x"{code[0x00002127-0x00002124,1]}", -- 0x00002124
    x"{code[0x0000212b-0x00002128,1]}", -- 0x00002128
    x"{code[0x0000212f-0x0000212c,1]}", -- 0x0000212c
    x"{code[0x00002133-0x00002130,1]}", -- 0x00002130
    x"{code[0x00002137-0x00002134,1]}", -- 0x00002134
    x"{code[0x0000213b-0x00002138,1]}", -- 0x00002138
    x"{code[0x0000213f-0x0000213c,1]}", -- 0x0000213c
    x"{code[0x00002143-0x00002140,1]}", -- 0x00002140
    x"{code[0x00002147-0x00002144,1]}", -- 0x00002144
    x"{code[0x0000214b-0x00002148,1]}", -- 0x00002148
    x"{code[0x0000214f-0x0000214c,1]}", -- 0x0000214c
    x"{code[0x00002153-0x00002150,1]}", -- 0x00002150
    x"{code[0x00002157-0x00002154,1]}", -- 0x00002154
    x"{code[0x0000215b-0x00002158,1]}", -- 0x00002158
    x"{code[0x0000215f-0x0000215c,1]}", -- 0x0000215c
    x"{code[0x00002163-0x00002160,1]}", -- 0x00002160
    x"{code[0x00002167-0x00002164,1]}", -- 0x00002164
    x"{code[0x0000216b-0x00002168,1]}", -- 0x00002168
    x"{code[0x0000216f-0x0000216c,1]}", -- 0x0000216c
    x"{code[0x00002173-0x00002170,1]}", -- 0x00002170
    x"{code[0x00002177-0x00002174,1]}", -- 0x00002174
    x"{code[0x0000217b-0x00002178,1]}", -- 0x00002178
    x"{code[0x0000217f-0x0000217c,1]}", -- 0x0000217c
    x"{code[0x00002183-0x00002180,1]}", -- 0x00002180
    x"{code[0x00002187-0x00002184,1]}", -- 0x00002184
    x"{code[0x0000218b-0x00002188,1]}", -- 0x00002188
    x"{code[0x0000218f-0x0000218c,1]}", -- 0x0000218c
    x"{code[0x00002193-0x00002190,1]}", -- 0x00002190
    x"{code[0x00002197-0x00002194,1]}", -- 0x00002194
    x"{code[0x0000219b-0x00002198,1]}", -- 0x00002198
    x"{code[0x0000219f-0x0000219c,1]}", -- 0x0000219c
    x"{code[0x000021a3-0x000021a0,1]}", -- 0x000021a0
    x"{code[0x000021a7-0x000021a4,1]}", -- 0x000021a4
    x"{code[0x000021ab-0x000021a8,1]}", -- 0x000021a8
    x"{code[0x000021af-0x000021ac,1]}", -- 0x000021ac
    x"{code[0x000021b3-0x000021b0,1]}", -- 0x000021b0
    x"{code[0x000021b7-0x000021b4,1]}", -- 0x000021b4
    x"{code[0x000021bb-0x000021b8,1]}", -- 0x000021b8
    x"{code[0x000021bf-0x000021bc,1]}", -- 0x000021bc
    x"{code[0x000021c3-0x000021c0,1]}", -- 0x000021c0
    x"{code[0x000021c7-0x000021c4,1]}", -- 0x000021c4
    x"{code[0x000021cb-0x000021c8,1]}", -- 0x000021c8
    x"{code[0x000021cf-0x000021cc,1]}", -- 0x000021cc
    x"{code[0x000021d3-0x000021d0,1]}", -- 0x000021d0
    x"{code[0x000021d7-0x000021d4,1]}", -- 0x000021d4
    x"{code[0x000021db-0x000021d8,1]}", -- 0x000021d8
    x"{code[0x000021df-0x000021dc,1]}", -- 0x000021dc
    x"{code[0x000021e3-0x000021e0,1]}", -- 0x000021e0
    x"{code[0x000021e7-0x000021e4,1]}", -- 0x000021e4
    x"{code[0x000021eb-0x000021e8,1]}", -- 0x000021e8
    x"{code[0x000021ef-0x000021ec,1]}", -- 0x000021ec
    x"{code[0x000021f3-0x000021f0,1]}", -- 0x000021f0
    x"{code[0x000021f7-0x000021f4,1]}", -- 0x000021f4
    x"{code[0x000021fb-0x000021f8,1]}", -- 0x000021f8
    x"{code[0x000021ff-0x000021fc,1]}", -- 0x000021fc
    x"{code[0x00002203-0x00002200,1]}", -- 0x00002200
    x"{code[0x00002207-0x00002204,1]}", -- 0x00002204
    x"{code[0x0000220b-0x00002208,1]}", -- 0x00002208
    x"{code[0x0000220f-0x0000220c,1]}", -- 0x0000220c
    x"{code[0x00002213-0x00002210,1]}", -- 0x00002210
    x"{code[0x00002217-0x00002214,1]}", -- 0x00002214
    x"{code[0x0000221b-0x00002218,1]}", -- 0x00002218
    x"{code[0x0000221f-0x0000221c,1]}", -- 0x0000221c
    x"{code[0x00002223-0x00002220,1]}", -- 0x00002220
    x"{code[0x00002227-0x00002224,1]}", -- 0x00002224
    x"{code[0x0000222b-0x00002228,1]}", -- 0x00002228
    x"{code[0x0000222f-0x0000222c,1]}", -- 0x0000222c
    x"{code[0x00002233-0x00002230,1]}", -- 0x00002230
    x"{code[0x00002237-0x00002234,1]}", -- 0x00002234
    x"{code[0x0000223b-0x00002238,1]}", -- 0x00002238
    x"{code[0x0000223f-0x0000223c,1]}", -- 0x0000223c
    x"{code[0x00002243-0x00002240,1]}", -- 0x00002240
    x"{code[0x00002247-0x00002244,1]}", -- 0x00002244
    x"{code[0x0000224b-0x00002248,1]}", -- 0x00002248
    x"{code[0x0000224f-0x0000224c,1]}", -- 0x0000224c
    x"{code[0x00002253-0x00002250,1]}", -- 0x00002250
    x"{code[0x00002257-0x00002254,1]}", -- 0x00002254
    x"{code[0x0000225b-0x00002258,1]}", -- 0x00002258
    x"{code[0x0000225f-0x0000225c,1]}", -- 0x0000225c
    x"{code[0x00002263-0x00002260,1]}", -- 0x00002260
    x"{code[0x00002267-0x00002264,1]}", -- 0x00002264
    x"{code[0x0000226b-0x00002268,1]}", -- 0x00002268
    x"{code[0x0000226f-0x0000226c,1]}", -- 0x0000226c
    x"{code[0x00002273-0x00002270,1]}", -- 0x00002270
    x"{code[0x00002277-0x00002274,1]}", -- 0x00002274
    x"{code[0x0000227b-0x00002278,1]}", -- 0x00002278
    x"{code[0x0000227f-0x0000227c,1]}", -- 0x0000227c
    x"{code[0x00002283-0x00002280,1]}", -- 0x00002280
    x"{code[0x00002287-0x00002284,1]}", -- 0x00002284
    x"{code[0x0000228b-0x00002288,1]}", -- 0x00002288
    x"{code[0x0000228f-0x0000228c,1]}", -- 0x0000228c
    x"{code[0x00002293-0x00002290,1]}", -- 0x00002290
    x"{code[0x00002297-0x00002294,1]}", -- 0x00002294
    x"{code[0x0000229b-0x00002298,1]}", -- 0x00002298
    x"{code[0x0000229f-0x0000229c,1]}", -- 0x0000229c
    x"{code[0x000022a3-0x000022a0,1]}", -- 0x000022a0
    x"{code[0x000022a7-0x000022a4,1]}", -- 0x000022a4
    x"{code[0x000022ab-0x000022a8,1]}", -- 0x000022a8
    x"{code[0x000022af-0x000022ac,1]}", -- 0x000022ac
    x"{code[0x000022b3-0x000022b0,1]}", -- 0x000022b0
    x"{code[0x000022b7-0x000022b4,1]}", -- 0x000022b4
    x"{code[0x000022bb-0x000022b8,1]}", -- 0x000022b8
    x"{code[0x000022bf-0x000022bc,1]}", -- 0x000022bc
    x"{code[0x000022c3-0x000022c0,1]}", -- 0x000022c0
    x"{code[0x000022c7-0x000022c4,1]}", -- 0x000022c4
    x"{code[0x000022cb-0x000022c8,1]}", -- 0x000022c8
    x"{code[0x000022cf-0x000022cc,1]}", -- 0x000022cc
    x"{code[0x000022d3-0x000022d0,1]}", -- 0x000022d0
    x"{code[0x000022d7-0x000022d4,1]}", -- 0x000022d4
    x"{code[0x000022db-0x000022d8,1]}", -- 0x000022d8
    x"{code[0x000022df-0x000022dc,1]}", -- 0x000022dc
    x"{code[0x000022e3-0x000022e0,1]}", -- 0x000022e0
    x"{code[0x000022e7-0x000022e4,1]}", -- 0x000022e4
    x"{code[0x000022eb-0x000022e8,1]}", -- 0x000022e8
    x"{code[0x000022ef-0x000022ec,1]}", -- 0x000022ec
    x"{code[0x000022f3-0x000022f0,1]}", -- 0x000022f0
    x"{code[0x000022f7-0x000022f4,1]}", -- 0x000022f4
    x"{code[0x000022fb-0x000022f8,1]}", -- 0x000022f8
    x"{code[0x000022ff-0x000022fc,1]}", -- 0x000022fc
    x"{code[0x00002303-0x00002300,1]}", -- 0x00002300
    x"{code[0x00002307-0x00002304,1]}", -- 0x00002304
    x"{code[0x0000230b-0x00002308,1]}", -- 0x00002308
    x"{code[0x0000230f-0x0000230c,1]}", -- 0x0000230c
    x"{code[0x00002313-0x00002310,1]}", -- 0x00002310
    x"{code[0x00002317-0x00002314,1]}", -- 0x00002314
    x"{code[0x0000231b-0x00002318,1]}", -- 0x00002318
    x"{code[0x0000231f-0x0000231c,1]}", -- 0x0000231c
    x"{code[0x00002323-0x00002320,1]}", -- 0x00002320
    x"{code[0x00002327-0x00002324,1]}", -- 0x00002324
    x"{code[0x0000232b-0x00002328,1]}", -- 0x00002328
    x"{code[0x0000232f-0x0000232c,1]}", -- 0x0000232c
    x"{code[0x00002333-0x00002330,1]}", -- 0x00002330
    x"{code[0x00002337-0x00002334,1]}", -- 0x00002334
    x"{code[0x0000233b-0x00002338,1]}", -- 0x00002338
    x"{code[0x0000233f-0x0000233c,1]}", -- 0x0000233c
    x"{code[0x00002343-0x00002340,1]}", -- 0x00002340
    x"{code[0x00002347-0x00002344,1]}", -- 0x00002344
    x"{code[0x0000234b-0x00002348,1]}", -- 0x00002348
    x"{code[0x0000234f-0x0000234c,1]}", -- 0x0000234c
    x"{code[0x00002353-0x00002350,1]}", -- 0x00002350
    x"{code[0x00002357-0x00002354,1]}", -- 0x00002354
    x"{code[0x0000235b-0x00002358,1]}", -- 0x00002358
    x"{code[0x0000235f-0x0000235c,1]}", -- 0x0000235c
    x"{code[0x00002363-0x00002360,1]}", -- 0x00002360
    x"{code[0x00002367-0x00002364,1]}", -- 0x00002364
    x"{code[0x0000236b-0x00002368,1]}", -- 0x00002368
    x"{code[0x0000236f-0x0000236c,1]}", -- 0x0000236c
    x"{code[0x00002373-0x00002370,1]}", -- 0x00002370
    x"{code[0x00002377-0x00002374,1]}", -- 0x00002374
    x"{code[0x0000237b-0x00002378,1]}", -- 0x00002378
    x"{code[0x0000237f-0x0000237c,1]}", -- 0x0000237c
    x"{code[0x00002383-0x00002380,1]}", -- 0x00002380
    x"{code[0x00002387-0x00002384,1]}", -- 0x00002384
    x"{code[0x0000238b-0x00002388,1]}", -- 0x00002388
    x"{code[0x0000238f-0x0000238c,1]}", -- 0x0000238c
    x"{code[0x00002393-0x00002390,1]}", -- 0x00002390
    x"{code[0x00002397-0x00002394,1]}", -- 0x00002394
    x"{code[0x0000239b-0x00002398,1]}", -- 0x00002398
    x"{code[0x0000239f-0x0000239c,1]}", -- 0x0000239c
    x"{code[0x000023a3-0x000023a0,1]}", -- 0x000023a0
    x"{code[0x000023a7-0x000023a4,1]}", -- 0x000023a4
    x"{code[0x000023ab-0x000023a8,1]}", -- 0x000023a8
    x"{code[0x000023af-0x000023ac,1]}", -- 0x000023ac
    x"{code[0x000023b3-0x000023b0,1]}", -- 0x000023b0
    x"{code[0x000023b7-0x000023b4,1]}", -- 0x000023b4
    x"{code[0x000023bb-0x000023b8,1]}", -- 0x000023b8
    x"{code[0x000023bf-0x000023bc,1]}", -- 0x000023bc
    x"{code[0x000023c3-0x000023c0,1]}", -- 0x000023c0
    x"{code[0x000023c7-0x000023c4,1]}", -- 0x000023c4
    x"{code[0x000023cb-0x000023c8,1]}", -- 0x000023c8
    x"{code[0x000023cf-0x000023cc,1]}", -- 0x000023cc
    x"{code[0x000023d3-0x000023d0,1]}", -- 0x000023d0
    x"{code[0x000023d7-0x000023d4,1]}", -- 0x000023d4
    x"{code[0x000023db-0x000023d8,1]}", -- 0x000023d8
    x"{code[0x000023df-0x000023dc,1]}", -- 0x000023dc
    x"{code[0x000023e3-0x000023e0,1]}", -- 0x000023e0
    x"{code[0x000023e7-0x000023e4,1]}", -- 0x000023e4
    x"{code[0x000023eb-0x000023e8,1]}", -- 0x000023e8
    x"{code[0x000023ef-0x000023ec,1]}", -- 0x000023ec
    x"{code[0x000023f3-0x000023f0,1]}", -- 0x000023f0
    x"{code[0x000023f7-0x000023f4,1]}", -- 0x000023f4
    x"{code[0x000023fb-0x000023f8,1]}", -- 0x000023f8
    x"{code[0x000023ff-0x000023fc,1]}", -- 0x000023fc
    x"{code[0x00002403-0x00002400,1]}", -- 0x00002400
    x"{code[0x00002407-0x00002404,1]}", -- 0x00002404
    x"{code[0x0000240b-0x00002408,1]}", -- 0x00002408
    x"{code[0x0000240f-0x0000240c,1]}", -- 0x0000240c
    x"{code[0x00002413-0x00002410,1]}", -- 0x00002410
    x"{code[0x00002417-0x00002414,1]}", -- 0x00002414
    x"{code[0x0000241b-0x00002418,1]}", -- 0x00002418
    x"{code[0x0000241f-0x0000241c,1]}", -- 0x0000241c
    x"{code[0x00002423-0x00002420,1]}", -- 0x00002420
    x"{code[0x00002427-0x00002424,1]}", -- 0x00002424
    x"{code[0x0000242b-0x00002428,1]}", -- 0x00002428
    x"{code[0x0000242f-0x0000242c,1]}", -- 0x0000242c
    x"{code[0x00002433-0x00002430,1]}", -- 0x00002430
    x"{code[0x00002437-0x00002434,1]}", -- 0x00002434
    x"{code[0x0000243b-0x00002438,1]}", -- 0x00002438
    x"{code[0x0000243f-0x0000243c,1]}", -- 0x0000243c
    x"{code[0x00002443-0x00002440,1]}", -- 0x00002440
    x"{code[0x00002447-0x00002444,1]}", -- 0x00002444
    x"{code[0x0000244b-0x00002448,1]}", -- 0x00002448
    x"{code[0x0000244f-0x0000244c,1]}", -- 0x0000244c
    x"{code[0x00002453-0x00002450,1]}", -- 0x00002450
    x"{code[0x00002457-0x00002454,1]}", -- 0x00002454
    x"{code[0x0000245b-0x00002458,1]}", -- 0x00002458
    x"{code[0x0000245f-0x0000245c,1]}", -- 0x0000245c
    x"{code[0x00002463-0x00002460,1]}", -- 0x00002460
    x"{code[0x00002467-0x00002464,1]}", -- 0x00002464
    x"{code[0x0000246b-0x00002468,1]}", -- 0x00002468
    x"{code[0x0000246f-0x0000246c,1]}", -- 0x0000246c
    x"{code[0x00002473-0x00002470,1]}", -- 0x00002470
    x"{code[0x00002477-0x00002474,1]}", -- 0x00002474
    x"{code[0x0000247b-0x00002478,1]}", -- 0x00002478
    x"{code[0x0000247f-0x0000247c,1]}", -- 0x0000247c
    x"{code[0x00002483-0x00002480,1]}", -- 0x00002480
    x"{code[0x00002487-0x00002484,1]}", -- 0x00002484
    x"{code[0x0000248b-0x00002488,1]}", -- 0x00002488
    x"{code[0x0000248f-0x0000248c,1]}", -- 0x0000248c
    x"{code[0x00002493-0x00002490,1]}", -- 0x00002490
    x"{code[0x00002497-0x00002494,1]}", -- 0x00002494
    x"{code[0x0000249b-0x00002498,1]}", -- 0x00002498
    x"{code[0x0000249f-0x0000249c,1]}", -- 0x0000249c
    x"{code[0x000024a3-0x000024a0,1]}", -- 0x000024a0
    x"{code[0x000024a7-0x000024a4,1]}", -- 0x000024a4
    x"{code[0x000024ab-0x000024a8,1]}", -- 0x000024a8
    x"{code[0x000024af-0x000024ac,1]}", -- 0x000024ac
    x"{code[0x000024b3-0x000024b0,1]}", -- 0x000024b0
    x"{code[0x000024b7-0x000024b4,1]}", -- 0x000024b4
    x"{code[0x000024bb-0x000024b8,1]}", -- 0x000024b8
    x"{code[0x000024bf-0x000024bc,1]}", -- 0x000024bc
    x"{code[0x000024c3-0x000024c0,1]}", -- 0x000024c0
    x"{code[0x000024c7-0x000024c4,1]}", -- 0x000024c4
    x"{code[0x000024cb-0x000024c8,1]}", -- 0x000024c8
    x"{code[0x000024cf-0x000024cc,1]}", -- 0x000024cc
    x"{code[0x000024d3-0x000024d0,1]}", -- 0x000024d0
    x"{code[0x000024d7-0x000024d4,1]}", -- 0x000024d4
    x"{code[0x000024db-0x000024d8,1]}", -- 0x000024d8
    x"{code[0x000024df-0x000024dc,1]}", -- 0x000024dc
    x"{code[0x000024e3-0x000024e0,1]}", -- 0x000024e0
    x"{code[0x000024e7-0x000024e4,1]}", -- 0x000024e4
    x"{code[0x000024eb-0x000024e8,1]}", -- 0x000024e8
    x"{code[0x000024ef-0x000024ec,1]}", -- 0x000024ec
    x"{code[0x000024f3-0x000024f0,1]}", -- 0x000024f0
    x"{code[0x000024f7-0x000024f4,1]}", -- 0x000024f4
    x"{code[0x000024fb-0x000024f8,1]}", -- 0x000024f8
    x"{code[0x000024ff-0x000024fc,1]}", -- 0x000024fc
    x"{code[0x00002503-0x00002500,1]}", -- 0x00002500
    x"{code[0x00002507-0x00002504,1]}", -- 0x00002504
    x"{code[0x0000250b-0x00002508,1]}", -- 0x00002508
    x"{code[0x0000250f-0x0000250c,1]}", -- 0x0000250c
    x"{code[0x00002513-0x00002510,1]}", -- 0x00002510
    x"{code[0x00002517-0x00002514,1]}", -- 0x00002514
    x"{code[0x0000251b-0x00002518,1]}", -- 0x00002518
    x"{code[0x0000251f-0x0000251c,1]}", -- 0x0000251c
    x"{code[0x00002523-0x00002520,1]}", -- 0x00002520
    x"{code[0x00002527-0x00002524,1]}", -- 0x00002524
    x"{code[0x0000252b-0x00002528,1]}", -- 0x00002528
    x"{code[0x0000252f-0x0000252c,1]}", -- 0x0000252c
    x"{code[0x00002533-0x00002530,1]}", -- 0x00002530
    x"{code[0x00002537-0x00002534,1]}", -- 0x00002534
    x"{code[0x0000253b-0x00002538,1]}", -- 0x00002538
    x"{code[0x0000253f-0x0000253c,1]}", -- 0x0000253c
    x"{code[0x00002543-0x00002540,1]}", -- 0x00002540
    x"{code[0x00002547-0x00002544,1]}", -- 0x00002544
    x"{code[0x0000254b-0x00002548,1]}", -- 0x00002548
    x"{code[0x0000254f-0x0000254c,1]}", -- 0x0000254c
    x"{code[0x00002553-0x00002550,1]}", -- 0x00002550
    x"{code[0x00002557-0x00002554,1]}", -- 0x00002554
    x"{code[0x0000255b-0x00002558,1]}", -- 0x00002558
    x"{code[0x0000255f-0x0000255c,1]}", -- 0x0000255c
    x"{code[0x00002563-0x00002560,1]}", -- 0x00002560
    x"{code[0x00002567-0x00002564,1]}", -- 0x00002564
    x"{code[0x0000256b-0x00002568,1]}", -- 0x00002568
    x"{code[0x0000256f-0x0000256c,1]}", -- 0x0000256c
    x"{code[0x00002573-0x00002570,1]}", -- 0x00002570
    x"{code[0x00002577-0x00002574,1]}", -- 0x00002574
    x"{code[0x0000257b-0x00002578,1]}", -- 0x00002578
    x"{code[0x0000257f-0x0000257c,1]}", -- 0x0000257c
    x"{code[0x00002583-0x00002580,1]}", -- 0x00002580
    x"{code[0x00002587-0x00002584,1]}", -- 0x00002584
    x"{code[0x0000258b-0x00002588,1]}", -- 0x00002588
    x"{code[0x0000258f-0x0000258c,1]}", -- 0x0000258c
    x"{code[0x00002593-0x00002590,1]}", -- 0x00002590
    x"{code[0x00002597-0x00002594,1]}", -- 0x00002594
    x"{code[0x0000259b-0x00002598,1]}", -- 0x00002598
    x"{code[0x0000259f-0x0000259c,1]}", -- 0x0000259c
    x"{code[0x000025a3-0x000025a0,1]}", -- 0x000025a0
    x"{code[0x000025a7-0x000025a4,1]}", -- 0x000025a4
    x"{code[0x000025ab-0x000025a8,1]}", -- 0x000025a8
    x"{code[0x000025af-0x000025ac,1]}", -- 0x000025ac
    x"{code[0x000025b3-0x000025b0,1]}", -- 0x000025b0
    x"{code[0x000025b7-0x000025b4,1]}", -- 0x000025b4
    x"{code[0x000025bb-0x000025b8,1]}", -- 0x000025b8
    x"{code[0x000025bf-0x000025bc,1]}", -- 0x000025bc
    x"{code[0x000025c3-0x000025c0,1]}", -- 0x000025c0
    x"{code[0x000025c7-0x000025c4,1]}", -- 0x000025c4
    x"{code[0x000025cb-0x000025c8,1]}", -- 0x000025c8
    x"{code[0x000025cf-0x000025cc,1]}", -- 0x000025cc
    x"{code[0x000025d3-0x000025d0,1]}", -- 0x000025d0
    x"{code[0x000025d7-0x000025d4,1]}", -- 0x000025d4
    x"{code[0x000025db-0x000025d8,1]}", -- 0x000025d8
    x"{code[0x000025df-0x000025dc,1]}", -- 0x000025dc
    x"{code[0x000025e3-0x000025e0,1]}", -- 0x000025e0
    x"{code[0x000025e7-0x000025e4,1]}", -- 0x000025e4
    x"{code[0x000025eb-0x000025e8,1]}", -- 0x000025e8
    x"{code[0x000025ef-0x000025ec,1]}", -- 0x000025ec
    x"{code[0x000025f3-0x000025f0,1]}", -- 0x000025f0
    x"{code[0x000025f7-0x000025f4,1]}", -- 0x000025f4
    x"{code[0x000025fb-0x000025f8,1]}", -- 0x000025f8
    x"{code[0x000025ff-0x000025fc,1]}", -- 0x000025fc
    x"{code[0x00002603-0x00002600,1]}", -- 0x00002600
    x"{code[0x00002607-0x00002604,1]}", -- 0x00002604
    x"{code[0x0000260b-0x00002608,1]}", -- 0x00002608
    x"{code[0x0000260f-0x0000260c,1]}", -- 0x0000260c
    x"{code[0x00002613-0x00002610,1]}", -- 0x00002610
    x"{code[0x00002617-0x00002614,1]}", -- 0x00002614
    x"{code[0x0000261b-0x00002618,1]}", -- 0x00002618
    x"{code[0x0000261f-0x0000261c,1]}", -- 0x0000261c
    x"{code[0x00002623-0x00002620,1]}", -- 0x00002620
    x"{code[0x00002627-0x00002624,1]}", -- 0x00002624
    x"{code[0x0000262b-0x00002628,1]}", -- 0x00002628
    x"{code[0x0000262f-0x0000262c,1]}", -- 0x0000262c
    x"{code[0x00002633-0x00002630,1]}", -- 0x00002630
    x"{code[0x00002637-0x00002634,1]}", -- 0x00002634
    x"{code[0x0000263b-0x00002638,1]}", -- 0x00002638
    x"{code[0x0000263f-0x0000263c,1]}", -- 0x0000263c
    x"{code[0x00002643-0x00002640,1]}", -- 0x00002640
    x"{code[0x00002647-0x00002644,1]}", -- 0x00002644
    x"{code[0x0000264b-0x00002648,1]}", -- 0x00002648
    x"{code[0x0000264f-0x0000264c,1]}", -- 0x0000264c
    x"{code[0x00002653-0x00002650,1]}", -- 0x00002650
    x"{code[0x00002657-0x00002654,1]}", -- 0x00002654
    x"{code[0x0000265b-0x00002658,1]}", -- 0x00002658
    x"{code[0x0000265f-0x0000265c,1]}", -- 0x0000265c
    x"{code[0x00002663-0x00002660,1]}", -- 0x00002660
    x"{code[0x00002667-0x00002664,1]}", -- 0x00002664
    x"{code[0x0000266b-0x00002668,1]}", -- 0x00002668
    x"{code[0x0000266f-0x0000266c,1]}", -- 0x0000266c
    x"{code[0x00002673-0x00002670,1]}", -- 0x00002670
    x"{code[0x00002677-0x00002674,1]}", -- 0x00002674
    x"{code[0x0000267b-0x00002678,1]}", -- 0x00002678
    x"{code[0x0000267f-0x0000267c,1]}", -- 0x0000267c
    x"{code[0x00002683-0x00002680,1]}", -- 0x00002680
    x"{code[0x00002687-0x00002684,1]}", -- 0x00002684
    x"{code[0x0000268b-0x00002688,1]}", -- 0x00002688
    x"{code[0x0000268f-0x0000268c,1]}", -- 0x0000268c
    x"{code[0x00002693-0x00002690,1]}", -- 0x00002690
    x"{code[0x00002697-0x00002694,1]}", -- 0x00002694
    x"{code[0x0000269b-0x00002698,1]}", -- 0x00002698
    x"{code[0x0000269f-0x0000269c,1]}", -- 0x0000269c
    x"{code[0x000026a3-0x000026a0,1]}", -- 0x000026a0
    x"{code[0x000026a7-0x000026a4,1]}", -- 0x000026a4
    x"{code[0x000026ab-0x000026a8,1]}", -- 0x000026a8
    x"{code[0x000026af-0x000026ac,1]}", -- 0x000026ac
    x"{code[0x000026b3-0x000026b0,1]}", -- 0x000026b0
    x"{code[0x000026b7-0x000026b4,1]}", -- 0x000026b4
    x"{code[0x000026bb-0x000026b8,1]}", -- 0x000026b8
    x"{code[0x000026bf-0x000026bc,1]}", -- 0x000026bc
    x"{code[0x000026c3-0x000026c0,1]}", -- 0x000026c0
    x"{code[0x000026c7-0x000026c4,1]}", -- 0x000026c4
    x"{code[0x000026cb-0x000026c8,1]}", -- 0x000026c8
    x"{code[0x000026cf-0x000026cc,1]}", -- 0x000026cc
    x"{code[0x000026d3-0x000026d0,1]}", -- 0x000026d0
    x"{code[0x000026d7-0x000026d4,1]}", -- 0x000026d4
    x"{code[0x000026db-0x000026d8,1]}", -- 0x000026d8
    x"{code[0x000026df-0x000026dc,1]}", -- 0x000026dc
    x"{code[0x000026e3-0x000026e0,1]}", -- 0x000026e0
    x"{code[0x000026e7-0x000026e4,1]}", -- 0x000026e4
    x"{code[0x000026eb-0x000026e8,1]}", -- 0x000026e8
    x"{code[0x000026ef-0x000026ec,1]}", -- 0x000026ec
    x"{code[0x000026f3-0x000026f0,1]}", -- 0x000026f0
    x"{code[0x000026f7-0x000026f4,1]}", -- 0x000026f4
    x"{code[0x000026fb-0x000026f8,1]}", -- 0x000026f8
    x"{code[0x000026ff-0x000026fc,1]}", -- 0x000026fc
    x"{code[0x00002703-0x00002700,1]}", -- 0x00002700
    x"{code[0x00002707-0x00002704,1]}", -- 0x00002704
    x"{code[0x0000270b-0x00002708,1]}", -- 0x00002708
    x"{code[0x0000270f-0x0000270c,1]}", -- 0x0000270c
    x"{code[0x00002713-0x00002710,1]}", -- 0x00002710
    x"{code[0x00002717-0x00002714,1]}", -- 0x00002714
    x"{code[0x0000271b-0x00002718,1]}", -- 0x00002718
    x"{code[0x0000271f-0x0000271c,1]}", -- 0x0000271c
    x"{code[0x00002723-0x00002720,1]}", -- 0x00002720
    x"{code[0x00002727-0x00002724,1]}", -- 0x00002724
    x"{code[0x0000272b-0x00002728,1]}", -- 0x00002728
    x"{code[0x0000272f-0x0000272c,1]}", -- 0x0000272c
    x"{code[0x00002733-0x00002730,1]}", -- 0x00002730
    x"{code[0x00002737-0x00002734,1]}", -- 0x00002734
    x"{code[0x0000273b-0x00002738,1]}", -- 0x00002738
    x"{code[0x0000273f-0x0000273c,1]}", -- 0x0000273c
    x"{code[0x00002743-0x00002740,1]}", -- 0x00002740
    x"{code[0x00002747-0x00002744,1]}", -- 0x00002744
    x"{code[0x0000274b-0x00002748,1]}", -- 0x00002748
    x"{code[0x0000274f-0x0000274c,1]}", -- 0x0000274c
    x"{code[0x00002753-0x00002750,1]}", -- 0x00002750
    x"{code[0x00002757-0x00002754,1]}", -- 0x00002754
    x"{code[0x0000275b-0x00002758,1]}", -- 0x00002758
    x"{code[0x0000275f-0x0000275c,1]}", -- 0x0000275c
    x"{code[0x00002763-0x00002760,1]}", -- 0x00002760
    x"{code[0x00002767-0x00002764,1]}", -- 0x00002764
    x"{code[0x0000276b-0x00002768,1]}", -- 0x00002768
    x"{code[0x0000276f-0x0000276c,1]}", -- 0x0000276c
    x"{code[0x00002773-0x00002770,1]}", -- 0x00002770
    x"{code[0x00002777-0x00002774,1]}", -- 0x00002774
    x"{code[0x0000277b-0x00002778,1]}", -- 0x00002778
    x"{code[0x0000277f-0x0000277c,1]}", -- 0x0000277c
    x"{code[0x00002783-0x00002780,1]}", -- 0x00002780
    x"{code[0x00002787-0x00002784,1]}", -- 0x00002784
    x"{code[0x0000278b-0x00002788,1]}", -- 0x00002788
    x"{code[0x0000278f-0x0000278c,1]}", -- 0x0000278c
    x"{code[0x00002793-0x00002790,1]}", -- 0x00002790
    x"{code[0x00002797-0x00002794,1]}", -- 0x00002794
    x"{code[0x0000279b-0x00002798,1]}", -- 0x00002798
    x"{code[0x0000279f-0x0000279c,1]}", -- 0x0000279c
    x"{code[0x000027a3-0x000027a0,1]}", -- 0x000027a0
    x"{code[0x000027a7-0x000027a4,1]}", -- 0x000027a4
    x"{code[0x000027ab-0x000027a8,1]}", -- 0x000027a8
    x"{code[0x000027af-0x000027ac,1]}", -- 0x000027ac
    x"{code[0x000027b3-0x000027b0,1]}", -- 0x000027b0
    x"{code[0x000027b7-0x000027b4,1]}", -- 0x000027b4
    x"{code[0x000027bb-0x000027b8,1]}", -- 0x000027b8
    x"{code[0x000027bf-0x000027bc,1]}", -- 0x000027bc
    x"{code[0x000027c3-0x000027c0,1]}", -- 0x000027c0
    x"{code[0x000027c7-0x000027c4,1]}", -- 0x000027c4
    x"{code[0x000027cb-0x000027c8,1]}", -- 0x000027c8
    x"{code[0x000027cf-0x000027cc,1]}", -- 0x000027cc
    x"{code[0x000027d3-0x000027d0,1]}", -- 0x000027d0
    x"{code[0x000027d7-0x000027d4,1]}", -- 0x000027d4
    x"{code[0x000027db-0x000027d8,1]}", -- 0x000027d8
    x"{code[0x000027df-0x000027dc,1]}", -- 0x000027dc
    x"{code[0x000027e3-0x000027e0,1]}", -- 0x000027e0
    x"{code[0x000027e7-0x000027e4,1]}", -- 0x000027e4
    x"{code[0x000027eb-0x000027e8,1]}", -- 0x000027e8
    x"{code[0x000027ef-0x000027ec,1]}", -- 0x000027ec
    x"{code[0x000027f3-0x000027f0,1]}", -- 0x000027f0
    x"{code[0x000027f7-0x000027f4,1]}", -- 0x000027f4
    x"{code[0x000027fb-0x000027f8,1]}", -- 0x000027f8
    x"{code[0x000027ff-0x000027fc,1]}", -- 0x000027fc
    x"{code[0x00002803-0x00002800,1]}", -- 0x00002800
    x"{code[0x00002807-0x00002804,1]}", -- 0x00002804
    x"{code[0x0000280b-0x00002808,1]}", -- 0x00002808
    x"{code[0x0000280f-0x0000280c,1]}", -- 0x0000280c
    x"{code[0x00002813-0x00002810,1]}", -- 0x00002810
    x"{code[0x00002817-0x00002814,1]}", -- 0x00002814
    x"{code[0x0000281b-0x00002818,1]}", -- 0x00002818
    x"{code[0x0000281f-0x0000281c,1]}", -- 0x0000281c
    x"{code[0x00002823-0x00002820,1]}", -- 0x00002820
    x"{code[0x00002827-0x00002824,1]}", -- 0x00002824
    x"{code[0x0000282b-0x00002828,1]}", -- 0x00002828
    x"{code[0x0000282f-0x0000282c,1]}", -- 0x0000282c
    x"{code[0x00002833-0x00002830,1]}", -- 0x00002830
    x"{code[0x00002837-0x00002834,1]}", -- 0x00002834
    x"{code[0x0000283b-0x00002838,1]}", -- 0x00002838
    x"{code[0x0000283f-0x0000283c,1]}", -- 0x0000283c
    x"{code[0x00002843-0x00002840,1]}", -- 0x00002840
    x"{code[0x00002847-0x00002844,1]}", -- 0x00002844
    x"{code[0x0000284b-0x00002848,1]}", -- 0x00002848
    x"{code[0x0000284f-0x0000284c,1]}", -- 0x0000284c
    x"{code[0x00002853-0x00002850,1]}", -- 0x00002850
    x"{code[0x00002857-0x00002854,1]}", -- 0x00002854
    x"{code[0x0000285b-0x00002858,1]}", -- 0x00002858
    x"{code[0x0000285f-0x0000285c,1]}", -- 0x0000285c
    x"{code[0x00002863-0x00002860,1]}", -- 0x00002860
    x"{code[0x00002867-0x00002864,1]}", -- 0x00002864
    x"{code[0x0000286b-0x00002868,1]}", -- 0x00002868
    x"{code[0x0000286f-0x0000286c,1]}", -- 0x0000286c
    x"{code[0x00002873-0x00002870,1]}", -- 0x00002870
    x"{code[0x00002877-0x00002874,1]}", -- 0x00002874
    x"{code[0x0000287b-0x00002878,1]}", -- 0x00002878
    x"{code[0x0000287f-0x0000287c,1]}", -- 0x0000287c
    x"{code[0x00002883-0x00002880,1]}", -- 0x00002880
    x"{code[0x00002887-0x00002884,1]}", -- 0x00002884
    x"{code[0x0000288b-0x00002888,1]}", -- 0x00002888
    x"{code[0x0000288f-0x0000288c,1]}", -- 0x0000288c
    x"{code[0x00002893-0x00002890,1]}", -- 0x00002890
    x"{code[0x00002897-0x00002894,1]}", -- 0x00002894
    x"{code[0x0000289b-0x00002898,1]}", -- 0x00002898
    x"{code[0x0000289f-0x0000289c,1]}", -- 0x0000289c
    x"{code[0x000028a3-0x000028a0,1]}", -- 0x000028a0
    x"{code[0x000028a7-0x000028a4,1]}", -- 0x000028a4
    x"{code[0x000028ab-0x000028a8,1]}", -- 0x000028a8
    x"{code[0x000028af-0x000028ac,1]}", -- 0x000028ac
    x"{code[0x000028b3-0x000028b0,1]}", -- 0x000028b0
    x"{code[0x000028b7-0x000028b4,1]}", -- 0x000028b4
    x"{code[0x000028bb-0x000028b8,1]}", -- 0x000028b8
    x"{code[0x000028bf-0x000028bc,1]}", -- 0x000028bc
    x"{code[0x000028c3-0x000028c0,1]}", -- 0x000028c0
    x"{code[0x000028c7-0x000028c4,1]}", -- 0x000028c4
    x"{code[0x000028cb-0x000028c8,1]}", -- 0x000028c8
    x"{code[0x000028cf-0x000028cc,1]}", -- 0x000028cc
    x"{code[0x000028d3-0x000028d0,1]}", -- 0x000028d0
    x"{code[0x000028d7-0x000028d4,1]}", -- 0x000028d4
    x"{code[0x000028db-0x000028d8,1]}", -- 0x000028d8
    x"{code[0x000028df-0x000028dc,1]}", -- 0x000028dc
    x"{code[0x000028e3-0x000028e0,1]}", -- 0x000028e0
    x"{code[0x000028e7-0x000028e4,1]}", -- 0x000028e4
    x"{code[0x000028eb-0x000028e8,1]}", -- 0x000028e8
    x"{code[0x000028ef-0x000028ec,1]}", -- 0x000028ec
    x"{code[0x000028f3-0x000028f0,1]}", -- 0x000028f0
    x"{code[0x000028f7-0x000028f4,1]}", -- 0x000028f4
    x"{code[0x000028fb-0x000028f8,1]}", -- 0x000028f8
    x"{code[0x000028ff-0x000028fc,1]}", -- 0x000028fc
    x"{code[0x00002903-0x00002900,1]}", -- 0x00002900
    x"{code[0x00002907-0x00002904,1]}", -- 0x00002904
    x"{code[0x0000290b-0x00002908,1]}", -- 0x00002908
    x"{code[0x0000290f-0x0000290c,1]}", -- 0x0000290c
    x"{code[0x00002913-0x00002910,1]}", -- 0x00002910
    x"{code[0x00002917-0x00002914,1]}", -- 0x00002914
    x"{code[0x0000291b-0x00002918,1]}", -- 0x00002918
    x"{code[0x0000291f-0x0000291c,1]}", -- 0x0000291c
    x"{code[0x00002923-0x00002920,1]}", -- 0x00002920
    x"{code[0x00002927-0x00002924,1]}", -- 0x00002924
    x"{code[0x0000292b-0x00002928,1]}", -- 0x00002928
    x"{code[0x0000292f-0x0000292c,1]}", -- 0x0000292c
    x"{code[0x00002933-0x00002930,1]}", -- 0x00002930
    x"{code[0x00002937-0x00002934,1]}", -- 0x00002934
    x"{code[0x0000293b-0x00002938,1]}", -- 0x00002938
    x"{code[0x0000293f-0x0000293c,1]}", -- 0x0000293c
    x"{code[0x00002943-0x00002940,1]}", -- 0x00002940
    x"{code[0x00002947-0x00002944,1]}", -- 0x00002944
    x"{code[0x0000294b-0x00002948,1]}", -- 0x00002948
    x"{code[0x0000294f-0x0000294c,1]}", -- 0x0000294c
    x"{code[0x00002953-0x00002950,1]}", -- 0x00002950
    x"{code[0x00002957-0x00002954,1]}", -- 0x00002954
    x"{code[0x0000295b-0x00002958,1]}", -- 0x00002958
    x"{code[0x0000295f-0x0000295c,1]}", -- 0x0000295c
    x"{code[0x00002963-0x00002960,1]}", -- 0x00002960
    x"{code[0x00002967-0x00002964,1]}", -- 0x00002964
    x"{code[0x0000296b-0x00002968,1]}", -- 0x00002968
    x"{code[0x0000296f-0x0000296c,1]}", -- 0x0000296c
    x"{code[0x00002973-0x00002970,1]}", -- 0x00002970
    x"{code[0x00002977-0x00002974,1]}", -- 0x00002974
    x"{code[0x0000297b-0x00002978,1]}", -- 0x00002978
    x"{code[0x0000297f-0x0000297c,1]}", -- 0x0000297c
    x"{code[0x00002983-0x00002980,1]}", -- 0x00002980
    x"{code[0x00002987-0x00002984,1]}", -- 0x00002984
    x"{code[0x0000298b-0x00002988,1]}", -- 0x00002988
    x"{code[0x0000298f-0x0000298c,1]}", -- 0x0000298c
    x"{code[0x00002993-0x00002990,1]}", -- 0x00002990
    x"{code[0x00002997-0x00002994,1]}", -- 0x00002994
    x"{code[0x0000299b-0x00002998,1]}", -- 0x00002998
    x"{code[0x0000299f-0x0000299c,1]}", -- 0x0000299c
    x"{code[0x000029a3-0x000029a0,1]}", -- 0x000029a0
    x"{code[0x000029a7-0x000029a4,1]}", -- 0x000029a4
    x"{code[0x000029ab-0x000029a8,1]}", -- 0x000029a8
    x"{code[0x000029af-0x000029ac,1]}", -- 0x000029ac
    x"{code[0x000029b3-0x000029b0,1]}", -- 0x000029b0
    x"{code[0x000029b7-0x000029b4,1]}", -- 0x000029b4
    x"{code[0x000029bb-0x000029b8,1]}", -- 0x000029b8
    x"{code[0x000029bf-0x000029bc,1]}", -- 0x000029bc
    x"{code[0x000029c3-0x000029c0,1]}", -- 0x000029c0
    x"{code[0x000029c7-0x000029c4,1]}", -- 0x000029c4
    x"{code[0x000029cb-0x000029c8,1]}", -- 0x000029c8
    x"{code[0x000029cf-0x000029cc,1]}", -- 0x000029cc
    x"{code[0x000029d3-0x000029d0,1]}", -- 0x000029d0
    x"{code[0x000029d7-0x000029d4,1]}", -- 0x000029d4
    x"{code[0x000029db-0x000029d8,1]}", -- 0x000029d8
    x"{code[0x000029df-0x000029dc,1]}", -- 0x000029dc
    x"{code[0x000029e3-0x000029e0,1]}", -- 0x000029e0
    x"{code[0x000029e7-0x000029e4,1]}", -- 0x000029e4
    x"{code[0x000029eb-0x000029e8,1]}", -- 0x000029e8
    x"{code[0x000029ef-0x000029ec,1]}", -- 0x000029ec
    x"{code[0x000029f3-0x000029f0,1]}", -- 0x000029f0
    x"{code[0x000029f7-0x000029f4,1]}", -- 0x000029f4
    x"{code[0x000029fb-0x000029f8,1]}", -- 0x000029f8
    x"{code[0x000029ff-0x000029fc,1]}", -- 0x000029fc
    x"{code[0x00002a03-0x00002a00,1]}", -- 0x00002a00
    x"{code[0x00002a07-0x00002a04,1]}", -- 0x00002a04
    x"{code[0x00002a0b-0x00002a08,1]}", -- 0x00002a08
    x"{code[0x00002a0f-0x00002a0c,1]}", -- 0x00002a0c
    x"{code[0x00002a13-0x00002a10,1]}", -- 0x00002a10
    x"{code[0x00002a17-0x00002a14,1]}", -- 0x00002a14
    x"{code[0x00002a1b-0x00002a18,1]}", -- 0x00002a18
    x"{code[0x00002a1f-0x00002a1c,1]}", -- 0x00002a1c
    x"{code[0x00002a23-0x00002a20,1]}", -- 0x00002a20
    x"{code[0x00002a27-0x00002a24,1]}", -- 0x00002a24
    x"{code[0x00002a2b-0x00002a28,1]}", -- 0x00002a28
    x"{code[0x00002a2f-0x00002a2c,1]}", -- 0x00002a2c
    x"{code[0x00002a33-0x00002a30,1]}", -- 0x00002a30
    x"{code[0x00002a37-0x00002a34,1]}", -- 0x00002a34
    x"{code[0x00002a3b-0x00002a38,1]}", -- 0x00002a38
    x"{code[0x00002a3f-0x00002a3c,1]}", -- 0x00002a3c
    x"{code[0x00002a43-0x00002a40,1]}", -- 0x00002a40
    x"{code[0x00002a47-0x00002a44,1]}", -- 0x00002a44
    x"{code[0x00002a4b-0x00002a48,1]}", -- 0x00002a48
    x"{code[0x00002a4f-0x00002a4c,1]}", -- 0x00002a4c
    x"{code[0x00002a53-0x00002a50,1]}", -- 0x00002a50
    x"{code[0x00002a57-0x00002a54,1]}", -- 0x00002a54
    x"{code[0x00002a5b-0x00002a58,1]}", -- 0x00002a58
    x"{code[0x00002a5f-0x00002a5c,1]}", -- 0x00002a5c
    x"{code[0x00002a63-0x00002a60,1]}", -- 0x00002a60
    x"{code[0x00002a67-0x00002a64,1]}", -- 0x00002a64
    x"{code[0x00002a6b-0x00002a68,1]}", -- 0x00002a68
    x"{code[0x00002a6f-0x00002a6c,1]}", -- 0x00002a6c
    x"{code[0x00002a73-0x00002a70,1]}", -- 0x00002a70
    x"{code[0x00002a77-0x00002a74,1]}", -- 0x00002a74
    x"{code[0x00002a7b-0x00002a78,1]}", -- 0x00002a78
    x"{code[0x00002a7f-0x00002a7c,1]}", -- 0x00002a7c
    x"{code[0x00002a83-0x00002a80,1]}", -- 0x00002a80
    x"{code[0x00002a87-0x00002a84,1]}", -- 0x00002a84
    x"{code[0x00002a8b-0x00002a88,1]}", -- 0x00002a88
    x"{code[0x00002a8f-0x00002a8c,1]}", -- 0x00002a8c
    x"{code[0x00002a93-0x00002a90,1]}", -- 0x00002a90
    x"{code[0x00002a97-0x00002a94,1]}", -- 0x00002a94
    x"{code[0x00002a9b-0x00002a98,1]}", -- 0x00002a98
    x"{code[0x00002a9f-0x00002a9c,1]}", -- 0x00002a9c
    x"{code[0x00002aa3-0x00002aa0,1]}", -- 0x00002aa0
    x"{code[0x00002aa7-0x00002aa4,1]}", -- 0x00002aa4
    x"{code[0x00002aab-0x00002aa8,1]}", -- 0x00002aa8
    x"{code[0x00002aaf-0x00002aac,1]}", -- 0x00002aac
    x"{code[0x00002ab3-0x00002ab0,1]}", -- 0x00002ab0
    x"{code[0x00002ab7-0x00002ab4,1]}", -- 0x00002ab4
    x"{code[0x00002abb-0x00002ab8,1]}", -- 0x00002ab8
    x"{code[0x00002abf-0x00002abc,1]}", -- 0x00002abc
    x"{code[0x00002ac3-0x00002ac0,1]}", -- 0x00002ac0
    x"{code[0x00002ac7-0x00002ac4,1]}", -- 0x00002ac4
    x"{code[0x00002acb-0x00002ac8,1]}", -- 0x00002ac8
    x"{code[0x00002acf-0x00002acc,1]}", -- 0x00002acc
    x"{code[0x00002ad3-0x00002ad0,1]}", -- 0x00002ad0
    x"{code[0x00002ad7-0x00002ad4,1]}", -- 0x00002ad4
    x"{code[0x00002adb-0x00002ad8,1]}", -- 0x00002ad8
    x"{code[0x00002adf-0x00002adc,1]}", -- 0x00002adc
    x"{code[0x00002ae3-0x00002ae0,1]}", -- 0x00002ae0
    x"{code[0x00002ae7-0x00002ae4,1]}", -- 0x00002ae4
    x"{code[0x00002aeb-0x00002ae8,1]}", -- 0x00002ae8
    x"{code[0x00002aef-0x00002aec,1]}", -- 0x00002aec
    x"{code[0x00002af3-0x00002af0,1]}", -- 0x00002af0
    x"{code[0x00002af7-0x00002af4,1]}", -- 0x00002af4
    x"{code[0x00002afb-0x00002af8,1]}", -- 0x00002af8
    x"{code[0x00002aff-0x00002afc,1]}", -- 0x00002afc
    x"{code[0x00002b03-0x00002b00,1]}", -- 0x00002b00
    x"{code[0x00002b07-0x00002b04,1]}", -- 0x00002b04
    x"{code[0x00002b0b-0x00002b08,1]}", -- 0x00002b08
    x"{code[0x00002b0f-0x00002b0c,1]}", -- 0x00002b0c
    x"{code[0x00002b13-0x00002b10,1]}", -- 0x00002b10
    x"{code[0x00002b17-0x00002b14,1]}", -- 0x00002b14
    x"{code[0x00002b1b-0x00002b18,1]}", -- 0x00002b18
    x"{code[0x00002b1f-0x00002b1c,1]}", -- 0x00002b1c
    x"{code[0x00002b23-0x00002b20,1]}", -- 0x00002b20
    x"{code[0x00002b27-0x00002b24,1]}", -- 0x00002b24
    x"{code[0x00002b2b-0x00002b28,1]}", -- 0x00002b28
    x"{code[0x00002b2f-0x00002b2c,1]}", -- 0x00002b2c
    x"{code[0x00002b33-0x00002b30,1]}", -- 0x00002b30
    x"{code[0x00002b37-0x00002b34,1]}", -- 0x00002b34
    x"{code[0x00002b3b-0x00002b38,1]}", -- 0x00002b38
    x"{code[0x00002b3f-0x00002b3c,1]}", -- 0x00002b3c
    x"{code[0x00002b43-0x00002b40,1]}", -- 0x00002b40
    x"{code[0x00002b47-0x00002b44,1]}", -- 0x00002b44
    x"{code[0x00002b4b-0x00002b48,1]}", -- 0x00002b48
    x"{code[0x00002b4f-0x00002b4c,1]}", -- 0x00002b4c
    x"{code[0x00002b53-0x00002b50,1]}", -- 0x00002b50
    x"{code[0x00002b57-0x00002b54,1]}", -- 0x00002b54
    x"{code[0x00002b5b-0x00002b58,1]}", -- 0x00002b58
    x"{code[0x00002b5f-0x00002b5c,1]}", -- 0x00002b5c
    x"{code[0x00002b63-0x00002b60,1]}", -- 0x00002b60
    x"{code[0x00002b67-0x00002b64,1]}", -- 0x00002b64
    x"{code[0x00002b6b-0x00002b68,1]}", -- 0x00002b68
    x"{code[0x00002b6f-0x00002b6c,1]}", -- 0x00002b6c
    x"{code[0x00002b73-0x00002b70,1]}", -- 0x00002b70
    x"{code[0x00002b77-0x00002b74,1]}", -- 0x00002b74
    x"{code[0x00002b7b-0x00002b78,1]}", -- 0x00002b78
    x"{code[0x00002b7f-0x00002b7c,1]}", -- 0x00002b7c
    x"{code[0x00002b83-0x00002b80,1]}", -- 0x00002b80
    x"{code[0x00002b87-0x00002b84,1]}", -- 0x00002b84
    x"{code[0x00002b8b-0x00002b88,1]}", -- 0x00002b88
    x"{code[0x00002b8f-0x00002b8c,1]}", -- 0x00002b8c
    x"{code[0x00002b93-0x00002b90,1]}", -- 0x00002b90
    x"{code[0x00002b97-0x00002b94,1]}", -- 0x00002b94
    x"{code[0x00002b9b-0x00002b98,1]}", -- 0x00002b98
    x"{code[0x00002b9f-0x00002b9c,1]}", -- 0x00002b9c
    x"{code[0x00002ba3-0x00002ba0,1]}", -- 0x00002ba0
    x"{code[0x00002ba7-0x00002ba4,1]}", -- 0x00002ba4
    x"{code[0x00002bab-0x00002ba8,1]}", -- 0x00002ba8
    x"{code[0x00002baf-0x00002bac,1]}", -- 0x00002bac
    x"{code[0x00002bb3-0x00002bb0,1]}", -- 0x00002bb0
    x"{code[0x00002bb7-0x00002bb4,1]}", -- 0x00002bb4
    x"{code[0x00002bbb-0x00002bb8,1]}", -- 0x00002bb8
    x"{code[0x00002bbf-0x00002bbc,1]}", -- 0x00002bbc
    x"{code[0x00002bc3-0x00002bc0,1]}", -- 0x00002bc0
    x"{code[0x00002bc7-0x00002bc4,1]}", -- 0x00002bc4
    x"{code[0x00002bcb-0x00002bc8,1]}", -- 0x00002bc8
    x"{code[0x00002bcf-0x00002bcc,1]}", -- 0x00002bcc
    x"{code[0x00002bd3-0x00002bd0,1]}", -- 0x00002bd0
    x"{code[0x00002bd7-0x00002bd4,1]}", -- 0x00002bd4
    x"{code[0x00002bdb-0x00002bd8,1]}", -- 0x00002bd8
    x"{code[0x00002bdf-0x00002bdc,1]}", -- 0x00002bdc
    x"{code[0x00002be3-0x00002be0,1]}", -- 0x00002be0
    x"{code[0x00002be7-0x00002be4,1]}", -- 0x00002be4
    x"{code[0x00002beb-0x00002be8,1]}", -- 0x00002be8
    x"{code[0x00002bef-0x00002bec,1]}", -- 0x00002bec
    x"{code[0x00002bf3-0x00002bf0,1]}", -- 0x00002bf0
    x"{code[0x00002bf7-0x00002bf4,1]}", -- 0x00002bf4
    x"{code[0x00002bfb-0x00002bf8,1]}", -- 0x00002bf8
    x"{code[0x00002bff-0x00002bfc,1]}", -- 0x00002bfc
    x"{code[0x00002c03-0x00002c00,1]}", -- 0x00002c00
    x"{code[0x00002c07-0x00002c04,1]}", -- 0x00002c04
    x"{code[0x00002c0b-0x00002c08,1]}", -- 0x00002c08
    x"{code[0x00002c0f-0x00002c0c,1]}", -- 0x00002c0c
    x"{code[0x00002c13-0x00002c10,1]}", -- 0x00002c10
    x"{code[0x00002c17-0x00002c14,1]}", -- 0x00002c14
    x"{code[0x00002c1b-0x00002c18,1]}", -- 0x00002c18
    x"{code[0x00002c1f-0x00002c1c,1]}", -- 0x00002c1c
    x"{code[0x00002c23-0x00002c20,1]}", -- 0x00002c20
    x"{code[0x00002c27-0x00002c24,1]}", -- 0x00002c24
    x"{code[0x00002c2b-0x00002c28,1]}", -- 0x00002c28
    x"{code[0x00002c2f-0x00002c2c,1]}", -- 0x00002c2c
    x"{code[0x00002c33-0x00002c30,1]}", -- 0x00002c30
    x"{code[0x00002c37-0x00002c34,1]}", -- 0x00002c34
    x"{code[0x00002c3b-0x00002c38,1]}", -- 0x00002c38
    x"{code[0x00002c3f-0x00002c3c,1]}", -- 0x00002c3c
    x"{code[0x00002c43-0x00002c40,1]}", -- 0x00002c40
    x"{code[0x00002c47-0x00002c44,1]}", -- 0x00002c44
    x"{code[0x00002c4b-0x00002c48,1]}", -- 0x00002c48
    x"{code[0x00002c4f-0x00002c4c,1]}", -- 0x00002c4c
    x"{code[0x00002c53-0x00002c50,1]}", -- 0x00002c50
    x"{code[0x00002c57-0x00002c54,1]}", -- 0x00002c54
    x"{code[0x00002c5b-0x00002c58,1]}", -- 0x00002c58
    x"{code[0x00002c5f-0x00002c5c,1]}", -- 0x00002c5c
    x"{code[0x00002c63-0x00002c60,1]}", -- 0x00002c60
    x"{code[0x00002c67-0x00002c64,1]}", -- 0x00002c64
    x"{code[0x00002c6b-0x00002c68,1]}", -- 0x00002c68
    x"{code[0x00002c6f-0x00002c6c,1]}", -- 0x00002c6c
    x"{code[0x00002c73-0x00002c70,1]}", -- 0x00002c70
    x"{code[0x00002c77-0x00002c74,1]}", -- 0x00002c74
    x"{code[0x00002c7b-0x00002c78,1]}", -- 0x00002c78
    x"{code[0x00002c7f-0x00002c7c,1]}", -- 0x00002c7c
    x"{code[0x00002c83-0x00002c80,1]}", -- 0x00002c80
    x"{code[0x00002c87-0x00002c84,1]}", -- 0x00002c84
    x"{code[0x00002c8b-0x00002c88,1]}", -- 0x00002c88
    x"{code[0x00002c8f-0x00002c8c,1]}", -- 0x00002c8c
    x"{code[0x00002c93-0x00002c90,1]}", -- 0x00002c90
    x"{code[0x00002c97-0x00002c94,1]}", -- 0x00002c94
    x"{code[0x00002c9b-0x00002c98,1]}", -- 0x00002c98
    x"{code[0x00002c9f-0x00002c9c,1]}", -- 0x00002c9c
    x"{code[0x00002ca3-0x00002ca0,1]}", -- 0x00002ca0
    x"{code[0x00002ca7-0x00002ca4,1]}", -- 0x00002ca4
    x"{code[0x00002cab-0x00002ca8,1]}", -- 0x00002ca8
    x"{code[0x00002caf-0x00002cac,1]}", -- 0x00002cac
    x"{code[0x00002cb3-0x00002cb0,1]}", -- 0x00002cb0
    x"{code[0x00002cb7-0x00002cb4,1]}", -- 0x00002cb4
    x"{code[0x00002cbb-0x00002cb8,1]}", -- 0x00002cb8
    x"{code[0x00002cbf-0x00002cbc,1]}", -- 0x00002cbc
    x"{code[0x00002cc3-0x00002cc0,1]}", -- 0x00002cc0
    x"{code[0x00002cc7-0x00002cc4,1]}", -- 0x00002cc4
    x"{code[0x00002ccb-0x00002cc8,1]}", -- 0x00002cc8
    x"{code[0x00002ccf-0x00002ccc,1]}", -- 0x00002ccc
    x"{code[0x00002cd3-0x00002cd0,1]}", -- 0x00002cd0
    x"{code[0x00002cd7-0x00002cd4,1]}", -- 0x00002cd4
    x"{code[0x00002cdb-0x00002cd8,1]}", -- 0x00002cd8
    x"{code[0x00002cdf-0x00002cdc,1]}", -- 0x00002cdc
    x"{code[0x00002ce3-0x00002ce0,1]}", -- 0x00002ce0
    x"{code[0x00002ce7-0x00002ce4,1]}", -- 0x00002ce4
    x"{code[0x00002ceb-0x00002ce8,1]}", -- 0x00002ce8
    x"{code[0x00002cef-0x00002cec,1]}", -- 0x00002cec
    x"{code[0x00002cf3-0x00002cf0,1]}", -- 0x00002cf0
    x"{code[0x00002cf7-0x00002cf4,1]}", -- 0x00002cf4
    x"{code[0x00002cfb-0x00002cf8,1]}", -- 0x00002cf8
    x"{code[0x00002cff-0x00002cfc,1]}", -- 0x00002cfc
    x"{code[0x00002d03-0x00002d00,1]}", -- 0x00002d00
    x"{code[0x00002d07-0x00002d04,1]}", -- 0x00002d04
    x"{code[0x00002d0b-0x00002d08,1]}", -- 0x00002d08
    x"{code[0x00002d0f-0x00002d0c,1]}", -- 0x00002d0c
    x"{code[0x00002d13-0x00002d10,1]}", -- 0x00002d10
    x"{code[0x00002d17-0x00002d14,1]}", -- 0x00002d14
    x"{code[0x00002d1b-0x00002d18,1]}", -- 0x00002d18
    x"{code[0x00002d1f-0x00002d1c,1]}", -- 0x00002d1c
    x"{code[0x00002d23-0x00002d20,1]}", -- 0x00002d20
    x"{code[0x00002d27-0x00002d24,1]}", -- 0x00002d24
    x"{code[0x00002d2b-0x00002d28,1]}", -- 0x00002d28
    x"{code[0x00002d2f-0x00002d2c,1]}", -- 0x00002d2c
    x"{code[0x00002d33-0x00002d30,1]}", -- 0x00002d30
    x"{code[0x00002d37-0x00002d34,1]}", -- 0x00002d34
    x"{code[0x00002d3b-0x00002d38,1]}", -- 0x00002d38
    x"{code[0x00002d3f-0x00002d3c,1]}", -- 0x00002d3c
    x"{code[0x00002d43-0x00002d40,1]}", -- 0x00002d40
    x"{code[0x00002d47-0x00002d44,1]}", -- 0x00002d44
    x"{code[0x00002d4b-0x00002d48,1]}", -- 0x00002d48
    x"{code[0x00002d4f-0x00002d4c,1]}", -- 0x00002d4c
    x"{code[0x00002d53-0x00002d50,1]}", -- 0x00002d50
    x"{code[0x00002d57-0x00002d54,1]}", -- 0x00002d54
    x"{code[0x00002d5b-0x00002d58,1]}", -- 0x00002d58
    x"{code[0x00002d5f-0x00002d5c,1]}", -- 0x00002d5c
    x"{code[0x00002d63-0x00002d60,1]}", -- 0x00002d60
    x"{code[0x00002d67-0x00002d64,1]}", -- 0x00002d64
    x"{code[0x00002d6b-0x00002d68,1]}", -- 0x00002d68
    x"{code[0x00002d6f-0x00002d6c,1]}", -- 0x00002d6c
    x"{code[0x00002d73-0x00002d70,1]}", -- 0x00002d70
    x"{code[0x00002d77-0x00002d74,1]}", -- 0x00002d74
    x"{code[0x00002d7b-0x00002d78,1]}", -- 0x00002d78
    x"{code[0x00002d7f-0x00002d7c,1]}", -- 0x00002d7c
    x"{code[0x00002d83-0x00002d80,1]}", -- 0x00002d80
    x"{code[0x00002d87-0x00002d84,1]}", -- 0x00002d84
    x"{code[0x00002d8b-0x00002d88,1]}", -- 0x00002d88
    x"{code[0x00002d8f-0x00002d8c,1]}", -- 0x00002d8c
    x"{code[0x00002d93-0x00002d90,1]}", -- 0x00002d90
    x"{code[0x00002d97-0x00002d94,1]}", -- 0x00002d94
    x"{code[0x00002d9b-0x00002d98,1]}", -- 0x00002d98
    x"{code[0x00002d9f-0x00002d9c,1]}", -- 0x00002d9c
    x"{code[0x00002da3-0x00002da0,1]}", -- 0x00002da0
    x"{code[0x00002da7-0x00002da4,1]}", -- 0x00002da4
    x"{code[0x00002dab-0x00002da8,1]}", -- 0x00002da8
    x"{code[0x00002daf-0x00002dac,1]}", -- 0x00002dac
    x"{code[0x00002db3-0x00002db0,1]}", -- 0x00002db0
    x"{code[0x00002db7-0x00002db4,1]}", -- 0x00002db4
    x"{code[0x00002dbb-0x00002db8,1]}", -- 0x00002db8
    x"{code[0x00002dbf-0x00002dbc,1]}", -- 0x00002dbc
    x"{code[0x00002dc3-0x00002dc0,1]}", -- 0x00002dc0
    x"{code[0x00002dc7-0x00002dc4,1]}", -- 0x00002dc4
    x"{code[0x00002dcb-0x00002dc8,1]}", -- 0x00002dc8
    x"{code[0x00002dcf-0x00002dcc,1]}", -- 0x00002dcc
    x"{code[0x00002dd3-0x00002dd0,1]}", -- 0x00002dd0
    x"{code[0x00002dd7-0x00002dd4,1]}", -- 0x00002dd4
    x"{code[0x00002ddb-0x00002dd8,1]}", -- 0x00002dd8
    x"{code[0x00002ddf-0x00002ddc,1]}", -- 0x00002ddc
    x"{code[0x00002de3-0x00002de0,1]}", -- 0x00002de0
    x"{code[0x00002de7-0x00002de4,1]}", -- 0x00002de4
    x"{code[0x00002deb-0x00002de8,1]}", -- 0x00002de8
    x"{code[0x00002def-0x00002dec,1]}", -- 0x00002dec
    x"{code[0x00002df3-0x00002df0,1]}", -- 0x00002df0
    x"{code[0x00002df7-0x00002df4,1]}", -- 0x00002df4
    x"{code[0x00002dfb-0x00002df8,1]}", -- 0x00002df8
    x"{code[0x00002dff-0x00002dfc,1]}", -- 0x00002dfc
    x"{code[0x00002e03-0x00002e00,1]}", -- 0x00002e00
    x"{code[0x00002e07-0x00002e04,1]}", -- 0x00002e04
    x"{code[0x00002e0b-0x00002e08,1]}", -- 0x00002e08
    x"{code[0x00002e0f-0x00002e0c,1]}", -- 0x00002e0c
    x"{code[0x00002e13-0x00002e10,1]}", -- 0x00002e10
    x"{code[0x00002e17-0x00002e14,1]}", -- 0x00002e14
    x"{code[0x00002e1b-0x00002e18,1]}", -- 0x00002e18
    x"{code[0x00002e1f-0x00002e1c,1]}", -- 0x00002e1c
    x"{code[0x00002e23-0x00002e20,1]}", -- 0x00002e20
    x"{code[0x00002e27-0x00002e24,1]}", -- 0x00002e24
    x"{code[0x00002e2b-0x00002e28,1]}", -- 0x00002e28
    x"{code[0x00002e2f-0x00002e2c,1]}", -- 0x00002e2c
    x"{code[0x00002e33-0x00002e30,1]}", -- 0x00002e30
    x"{code[0x00002e37-0x00002e34,1]}", -- 0x00002e34
    x"{code[0x00002e3b-0x00002e38,1]}", -- 0x00002e38
    x"{code[0x00002e3f-0x00002e3c,1]}", -- 0x00002e3c
    x"{code[0x00002e43-0x00002e40,1]}", -- 0x00002e40
    x"{code[0x00002e47-0x00002e44,1]}", -- 0x00002e44
    x"{code[0x00002e4b-0x00002e48,1]}", -- 0x00002e48
    x"{code[0x00002e4f-0x00002e4c,1]}", -- 0x00002e4c
    x"{code[0x00002e53-0x00002e50,1]}", -- 0x00002e50
    x"{code[0x00002e57-0x00002e54,1]}", -- 0x00002e54
    x"{code[0x00002e5b-0x00002e58,1]}", -- 0x00002e58
    x"{code[0x00002e5f-0x00002e5c,1]}", -- 0x00002e5c
    x"{code[0x00002e63-0x00002e60,1]}", -- 0x00002e60
    x"{code[0x00002e67-0x00002e64,1]}", -- 0x00002e64
    x"{code[0x00002e6b-0x00002e68,1]}", -- 0x00002e68
    x"{code[0x00002e6f-0x00002e6c,1]}", -- 0x00002e6c
    x"{code[0x00002e73-0x00002e70,1]}", -- 0x00002e70
    x"{code[0x00002e77-0x00002e74,1]}", -- 0x00002e74
    x"{code[0x00002e7b-0x00002e78,1]}", -- 0x00002e78
    x"{code[0x00002e7f-0x00002e7c,1]}", -- 0x00002e7c
    x"{code[0x00002e83-0x00002e80,1]}", -- 0x00002e80
    x"{code[0x00002e87-0x00002e84,1]}", -- 0x00002e84
    x"{code[0x00002e8b-0x00002e88,1]}", -- 0x00002e88
    x"{code[0x00002e8f-0x00002e8c,1]}", -- 0x00002e8c
    x"{code[0x00002e93-0x00002e90,1]}", -- 0x00002e90
    x"{code[0x00002e97-0x00002e94,1]}", -- 0x00002e94
    x"{code[0x00002e9b-0x00002e98,1]}", -- 0x00002e98
    x"{code[0x00002e9f-0x00002e9c,1]}", -- 0x00002e9c
    x"{code[0x00002ea3-0x00002ea0,1]}", -- 0x00002ea0
    x"{code[0x00002ea7-0x00002ea4,1]}", -- 0x00002ea4
    x"{code[0x00002eab-0x00002ea8,1]}", -- 0x00002ea8
    x"{code[0x00002eaf-0x00002eac,1]}", -- 0x00002eac
    x"{code[0x00002eb3-0x00002eb0,1]}", -- 0x00002eb0
    x"{code[0x00002eb7-0x00002eb4,1]}", -- 0x00002eb4
    x"{code[0x00002ebb-0x00002eb8,1]}", -- 0x00002eb8
    x"{code[0x00002ebf-0x00002ebc,1]}", -- 0x00002ebc
    x"{code[0x00002ec3-0x00002ec0,1]}", -- 0x00002ec0
    x"{code[0x00002ec7-0x00002ec4,1]}", -- 0x00002ec4
    x"{code[0x00002ecb-0x00002ec8,1]}", -- 0x00002ec8
    x"{code[0x00002ecf-0x00002ecc,1]}", -- 0x00002ecc
    x"{code[0x00002ed3-0x00002ed0,1]}", -- 0x00002ed0
    x"{code[0x00002ed7-0x00002ed4,1]}", -- 0x00002ed4
    x"{code[0x00002edb-0x00002ed8,1]}", -- 0x00002ed8
    x"{code[0x00002edf-0x00002edc,1]}", -- 0x00002edc
    x"{code[0x00002ee3-0x00002ee0,1]}", -- 0x00002ee0
    x"{code[0x00002ee7-0x00002ee4,1]}", -- 0x00002ee4
    x"{code[0x00002eeb-0x00002ee8,1]}", -- 0x00002ee8
    x"{code[0x00002eef-0x00002eec,1]}", -- 0x00002eec
    x"{code[0x00002ef3-0x00002ef0,1]}", -- 0x00002ef0
    x"{code[0x00002ef7-0x00002ef4,1]}", -- 0x00002ef4
    x"{code[0x00002efb-0x00002ef8,1]}", -- 0x00002ef8
    x"{code[0x00002eff-0x00002efc,1]}", -- 0x00002efc
    x"{code[0x00002f03-0x00002f00,1]}", -- 0x00002f00
    x"{code[0x00002f07-0x00002f04,1]}", -- 0x00002f04
    x"{code[0x00002f0b-0x00002f08,1]}", -- 0x00002f08
    x"{code[0x00002f0f-0x00002f0c,1]}", -- 0x00002f0c
    x"{code[0x00002f13-0x00002f10,1]}", -- 0x00002f10
    x"{code[0x00002f17-0x00002f14,1]}", -- 0x00002f14
    x"{code[0x00002f1b-0x00002f18,1]}", -- 0x00002f18
    x"{code[0x00002f1f-0x00002f1c,1]}", -- 0x00002f1c
    x"{code[0x00002f23-0x00002f20,1]}", -- 0x00002f20
    x"{code[0x00002f27-0x00002f24,1]}", -- 0x00002f24
    x"{code[0x00002f2b-0x00002f28,1]}", -- 0x00002f28
    x"{code[0x00002f2f-0x00002f2c,1]}", -- 0x00002f2c
    x"{code[0x00002f33-0x00002f30,1]}", -- 0x00002f30
    x"{code[0x00002f37-0x00002f34,1]}", -- 0x00002f34
    x"{code[0x00002f3b-0x00002f38,1]}", -- 0x00002f38
    x"{code[0x00002f3f-0x00002f3c,1]}", -- 0x00002f3c
    x"{code[0x00002f43-0x00002f40,1]}", -- 0x00002f40
    x"{code[0x00002f47-0x00002f44,1]}", -- 0x00002f44
    x"{code[0x00002f4b-0x00002f48,1]}", -- 0x00002f48
    x"{code[0x00002f4f-0x00002f4c,1]}", -- 0x00002f4c
    x"{code[0x00002f53-0x00002f50,1]}", -- 0x00002f50
    x"{code[0x00002f57-0x00002f54,1]}", -- 0x00002f54
    x"{code[0x00002f5b-0x00002f58,1]}", -- 0x00002f58
    x"{code[0x00002f5f-0x00002f5c,1]}", -- 0x00002f5c
    x"{code[0x00002f63-0x00002f60,1]}", -- 0x00002f60
    x"{code[0x00002f67-0x00002f64,1]}", -- 0x00002f64
    x"{code[0x00002f6b-0x00002f68,1]}", -- 0x00002f68
    x"{code[0x00002f6f-0x00002f6c,1]}", -- 0x00002f6c
    x"{code[0x00002f73-0x00002f70,1]}", -- 0x00002f70
    x"{code[0x00002f77-0x00002f74,1]}", -- 0x00002f74
    x"{code[0x00002f7b-0x00002f78,1]}", -- 0x00002f78
    x"{code[0x00002f7f-0x00002f7c,1]}", -- 0x00002f7c
    x"{code[0x00002f83-0x00002f80,1]}", -- 0x00002f80
    x"{code[0x00002f87-0x00002f84,1]}", -- 0x00002f84
    x"{code[0x00002f8b-0x00002f88,1]}", -- 0x00002f88
    x"{code[0x00002f8f-0x00002f8c,1]}", -- 0x00002f8c
    x"{code[0x00002f93-0x00002f90,1]}", -- 0x00002f90
    x"{code[0x00002f97-0x00002f94,1]}", -- 0x00002f94
    x"{code[0x00002f9b-0x00002f98,1]}", -- 0x00002f98
    x"{code[0x00002f9f-0x00002f9c,1]}", -- 0x00002f9c
    x"{code[0x00002fa3-0x00002fa0,1]}", -- 0x00002fa0
    x"{code[0x00002fa7-0x00002fa4,1]}", -- 0x00002fa4
    x"{code[0x00002fab-0x00002fa8,1]}", -- 0x00002fa8
    x"{code[0x00002faf-0x00002fac,1]}", -- 0x00002fac
    x"{code[0x00002fb3-0x00002fb0,1]}", -- 0x00002fb0
    x"{code[0x00002fb7-0x00002fb4,1]}", -- 0x00002fb4
    x"{code[0x00002fbb-0x00002fb8,1]}", -- 0x00002fb8
    x"{code[0x00002fbf-0x00002fbc,1]}", -- 0x00002fbc
    x"{code[0x00002fc3-0x00002fc0,1]}", -- 0x00002fc0
    x"{code[0x00002fc7-0x00002fc4,1]}", -- 0x00002fc4
    x"{code[0x00002fcb-0x00002fc8,1]}", -- 0x00002fc8
    x"{code[0x00002fcf-0x00002fcc,1]}", -- 0x00002fcc
    x"{code[0x00002fd3-0x00002fd0,1]}", -- 0x00002fd0
    x"{code[0x00002fd7-0x00002fd4,1]}", -- 0x00002fd4
    x"{code[0x00002fdb-0x00002fd8,1]}", -- 0x00002fd8
    x"{code[0x00002fdf-0x00002fdc,1]}", -- 0x00002fdc
    x"{code[0x00002fe3-0x00002fe0,1]}", -- 0x00002fe0
    x"{code[0x00002fe7-0x00002fe4,1]}", -- 0x00002fe4
    x"{code[0x00002feb-0x00002fe8,1]}", -- 0x00002fe8
    x"{code[0x00002fef-0x00002fec,1]}", -- 0x00002fec
    x"{code[0x00002ff3-0x00002ff0,1]}", -- 0x00002ff0
    x"{code[0x00002ff7-0x00002ff4,1]}", -- 0x00002ff4
    x"{code[0x00002ffb-0x00002ff8,1]}", -- 0x00002ff8
    x"{code[0x00002fff-0x00002ffc,1]}", -- 0x00002ffc
    x"{code[0x00003003-0x00003000,1]}", -- 0x00003000
    x"{code[0x00003007-0x00003004,1]}", -- 0x00003004
    x"{code[0x0000300b-0x00003008,1]}", -- 0x00003008
    x"{code[0x0000300f-0x0000300c,1]}", -- 0x0000300c
    x"{code[0x00003013-0x00003010,1]}", -- 0x00003010
    x"{code[0x00003017-0x00003014,1]}", -- 0x00003014
    x"{code[0x0000301b-0x00003018,1]}", -- 0x00003018
    x"{code[0x0000301f-0x0000301c,1]}", -- 0x0000301c
    x"{code[0x00003023-0x00003020,1]}", -- 0x00003020
    x"{code[0x00003027-0x00003024,1]}", -- 0x00003024
    x"{code[0x0000302b-0x00003028,1]}", -- 0x00003028
    x"{code[0x0000302f-0x0000302c,1]}", -- 0x0000302c
    x"{code[0x00003033-0x00003030,1]}", -- 0x00003030
    x"{code[0x00003037-0x00003034,1]}", -- 0x00003034
    x"{code[0x0000303b-0x00003038,1]}", -- 0x00003038
    x"{code[0x0000303f-0x0000303c,1]}", -- 0x0000303c
    x"{code[0x00003043-0x00003040,1]}", -- 0x00003040
    x"{code[0x00003047-0x00003044,1]}", -- 0x00003044
    x"{code[0x0000304b-0x00003048,1]}", -- 0x00003048
    x"{code[0x0000304f-0x0000304c,1]}", -- 0x0000304c
    x"{code[0x00003053-0x00003050,1]}", -- 0x00003050
    x"{code[0x00003057-0x00003054,1]}", -- 0x00003054
    x"{code[0x0000305b-0x00003058,1]}", -- 0x00003058
    x"{code[0x0000305f-0x0000305c,1]}", -- 0x0000305c
    x"{code[0x00003063-0x00003060,1]}", -- 0x00003060
    x"{code[0x00003067-0x00003064,1]}", -- 0x00003064
    x"{code[0x0000306b-0x00003068,1]}", -- 0x00003068
    x"{code[0x0000306f-0x0000306c,1]}", -- 0x0000306c
    x"{code[0x00003073-0x00003070,1]}", -- 0x00003070
    x"{code[0x00003077-0x00003074,1]}", -- 0x00003074
    x"{code[0x0000307b-0x00003078,1]}", -- 0x00003078
    x"{code[0x0000307f-0x0000307c,1]}", -- 0x0000307c
    x"{code[0x00003083-0x00003080,1]}", -- 0x00003080
    x"{code[0x00003087-0x00003084,1]}", -- 0x00003084
    x"{code[0x0000308b-0x00003088,1]}", -- 0x00003088
    x"{code[0x0000308f-0x0000308c,1]}", -- 0x0000308c
    x"{code[0x00003093-0x00003090,1]}", -- 0x00003090
    x"{code[0x00003097-0x00003094,1]}", -- 0x00003094
    x"{code[0x0000309b-0x00003098,1]}", -- 0x00003098
    x"{code[0x0000309f-0x0000309c,1]}", -- 0x0000309c
    x"{code[0x000030a3-0x000030a0,1]}", -- 0x000030a0
    x"{code[0x000030a7-0x000030a4,1]}", -- 0x000030a4
    x"{code[0x000030ab-0x000030a8,1]}", -- 0x000030a8
    x"{code[0x000030af-0x000030ac,1]}", -- 0x000030ac
    x"{code[0x000030b3-0x000030b0,1]}", -- 0x000030b0
    x"{code[0x000030b7-0x000030b4,1]}", -- 0x000030b4
    x"{code[0x000030bb-0x000030b8,1]}", -- 0x000030b8
    x"{code[0x000030bf-0x000030bc,1]}", -- 0x000030bc
    x"{code[0x000030c3-0x000030c0,1]}", -- 0x000030c0
    x"{code[0x000030c7-0x000030c4,1]}", -- 0x000030c4
    x"{code[0x000030cb-0x000030c8,1]}", -- 0x000030c8
    x"{code[0x000030cf-0x000030cc,1]}", -- 0x000030cc
    x"{code[0x000030d3-0x000030d0,1]}", -- 0x000030d0
    x"{code[0x000030d7-0x000030d4,1]}", -- 0x000030d4
    x"{code[0x000030db-0x000030d8,1]}", -- 0x000030d8
    x"{code[0x000030df-0x000030dc,1]}", -- 0x000030dc
    x"{code[0x000030e3-0x000030e0,1]}", -- 0x000030e0
    x"{code[0x000030e7-0x000030e4,1]}", -- 0x000030e4
    x"{code[0x000030eb-0x000030e8,1]}", -- 0x000030e8
    x"{code[0x000030ef-0x000030ec,1]}", -- 0x000030ec
    x"{code[0x000030f3-0x000030f0,1]}", -- 0x000030f0
    x"{code[0x000030f7-0x000030f4,1]}", -- 0x000030f4
    x"{code[0x000030fb-0x000030f8,1]}", -- 0x000030f8
    x"{code[0x000030ff-0x000030fc,1]}", -- 0x000030fc
    x"{code[0x00003103-0x00003100,1]}", -- 0x00003100
    x"{code[0x00003107-0x00003104,1]}", -- 0x00003104
    x"{code[0x0000310b-0x00003108,1]}", -- 0x00003108
    x"{code[0x0000310f-0x0000310c,1]}", -- 0x0000310c
    x"{code[0x00003113-0x00003110,1]}", -- 0x00003110
    x"{code[0x00003117-0x00003114,1]}", -- 0x00003114
    x"{code[0x0000311b-0x00003118,1]}", -- 0x00003118
    x"{code[0x0000311f-0x0000311c,1]}", -- 0x0000311c
    x"{code[0x00003123-0x00003120,1]}", -- 0x00003120
    x"{code[0x00003127-0x00003124,1]}", -- 0x00003124
    x"{code[0x0000312b-0x00003128,1]}", -- 0x00003128
    x"{code[0x0000312f-0x0000312c,1]}", -- 0x0000312c
    x"{code[0x00003133-0x00003130,1]}", -- 0x00003130
    x"{code[0x00003137-0x00003134,1]}", -- 0x00003134
    x"{code[0x0000313b-0x00003138,1]}", -- 0x00003138
    x"{code[0x0000313f-0x0000313c,1]}", -- 0x0000313c
    x"{code[0x00003143-0x00003140,1]}", -- 0x00003140
    x"{code[0x00003147-0x00003144,1]}", -- 0x00003144
    x"{code[0x0000314b-0x00003148,1]}", -- 0x00003148
    x"{code[0x0000314f-0x0000314c,1]}", -- 0x0000314c
    x"{code[0x00003153-0x00003150,1]}", -- 0x00003150
    x"{code[0x00003157-0x00003154,1]}", -- 0x00003154
    x"{code[0x0000315b-0x00003158,1]}", -- 0x00003158
    x"{code[0x0000315f-0x0000315c,1]}", -- 0x0000315c
    x"{code[0x00003163-0x00003160,1]}", -- 0x00003160
    x"{code[0x00003167-0x00003164,1]}", -- 0x00003164
    x"{code[0x0000316b-0x00003168,1]}", -- 0x00003168
    x"{code[0x0000316f-0x0000316c,1]}", -- 0x0000316c
    x"{code[0x00003173-0x00003170,1]}", -- 0x00003170
    x"{code[0x00003177-0x00003174,1]}", -- 0x00003174
    x"{code[0x0000317b-0x00003178,1]}", -- 0x00003178
    x"{code[0x0000317f-0x0000317c,1]}", -- 0x0000317c
    x"{code[0x00003183-0x00003180,1]}", -- 0x00003180
    x"{code[0x00003187-0x00003184,1]}", -- 0x00003184
    x"{code[0x0000318b-0x00003188,1]}", -- 0x00003188
    x"{code[0x0000318f-0x0000318c,1]}", -- 0x0000318c
    x"{code[0x00003193-0x00003190,1]}", -- 0x00003190
    x"{code[0x00003197-0x00003194,1]}", -- 0x00003194
    x"{code[0x0000319b-0x00003198,1]}", -- 0x00003198
    x"{code[0x0000319f-0x0000319c,1]}", -- 0x0000319c
    x"{code[0x000031a3-0x000031a0,1]}", -- 0x000031a0
    x"{code[0x000031a7-0x000031a4,1]}", -- 0x000031a4
    x"{code[0x000031ab-0x000031a8,1]}", -- 0x000031a8
    x"{code[0x000031af-0x000031ac,1]}", -- 0x000031ac
    x"{code[0x000031b3-0x000031b0,1]}", -- 0x000031b0
    x"{code[0x000031b7-0x000031b4,1]}", -- 0x000031b4
    x"{code[0x000031bb-0x000031b8,1]}", -- 0x000031b8
    x"{code[0x000031bf-0x000031bc,1]}", -- 0x000031bc
    x"{code[0x000031c3-0x000031c0,1]}", -- 0x000031c0
    x"{code[0x000031c7-0x000031c4,1]}", -- 0x000031c4
    x"{code[0x000031cb-0x000031c8,1]}", -- 0x000031c8
    x"{code[0x000031cf-0x000031cc,1]}", -- 0x000031cc
    x"{code[0x000031d3-0x000031d0,1]}", -- 0x000031d0
    x"{code[0x000031d7-0x000031d4,1]}", -- 0x000031d4
    x"{code[0x000031db-0x000031d8,1]}", -- 0x000031d8
    x"{code[0x000031df-0x000031dc,1]}", -- 0x000031dc
    x"{code[0x000031e3-0x000031e0,1]}", -- 0x000031e0
    x"{code[0x000031e7-0x000031e4,1]}", -- 0x000031e4
    x"{code[0x000031eb-0x000031e8,1]}", -- 0x000031e8
    x"{code[0x000031ef-0x000031ec,1]}", -- 0x000031ec
    x"{code[0x000031f3-0x000031f0,1]}", -- 0x000031f0
    x"{code[0x000031f7-0x000031f4,1]}", -- 0x000031f4
    x"{code[0x000031fb-0x000031f8,1]}", -- 0x000031f8
    x"{code[0x000031ff-0x000031fc,1]}", -- 0x000031fc
    x"{code[0x00003203-0x00003200,1]}", -- 0x00003200
    x"{code[0x00003207-0x00003204,1]}", -- 0x00003204
    x"{code[0x0000320b-0x00003208,1]}", -- 0x00003208
    x"{code[0x0000320f-0x0000320c,1]}", -- 0x0000320c
    x"{code[0x00003213-0x00003210,1]}", -- 0x00003210
    x"{code[0x00003217-0x00003214,1]}", -- 0x00003214
    x"{code[0x0000321b-0x00003218,1]}", -- 0x00003218
    x"{code[0x0000321f-0x0000321c,1]}", -- 0x0000321c
    x"{code[0x00003223-0x00003220,1]}", -- 0x00003220
    x"{code[0x00003227-0x00003224,1]}", -- 0x00003224
    x"{code[0x0000322b-0x00003228,1]}", -- 0x00003228
    x"{code[0x0000322f-0x0000322c,1]}", -- 0x0000322c
    x"{code[0x00003233-0x00003230,1]}", -- 0x00003230
    x"{code[0x00003237-0x00003234,1]}", -- 0x00003234
    x"{code[0x0000323b-0x00003238,1]}", -- 0x00003238
    x"{code[0x0000323f-0x0000323c,1]}", -- 0x0000323c
    x"{code[0x00003243-0x00003240,1]}", -- 0x00003240
    x"{code[0x00003247-0x00003244,1]}", -- 0x00003244
    x"{code[0x0000324b-0x00003248,1]}", -- 0x00003248
    x"{code[0x0000324f-0x0000324c,1]}", -- 0x0000324c
    x"{code[0x00003253-0x00003250,1]}", -- 0x00003250
    x"{code[0x00003257-0x00003254,1]}", -- 0x00003254
    x"{code[0x0000325b-0x00003258,1]}", -- 0x00003258
    x"{code[0x0000325f-0x0000325c,1]}", -- 0x0000325c
    x"{code[0x00003263-0x00003260,1]}", -- 0x00003260
    x"{code[0x00003267-0x00003264,1]}", -- 0x00003264
    x"{code[0x0000326b-0x00003268,1]}", -- 0x00003268
    x"{code[0x0000326f-0x0000326c,1]}", -- 0x0000326c
    x"{code[0x00003273-0x00003270,1]}", -- 0x00003270
    x"{code[0x00003277-0x00003274,1]}", -- 0x00003274
    x"{code[0x0000327b-0x00003278,1]}", -- 0x00003278
    x"{code[0x0000327f-0x0000327c,1]}", -- 0x0000327c
    x"{code[0x00003283-0x00003280,1]}", -- 0x00003280
    x"{code[0x00003287-0x00003284,1]}", -- 0x00003284
    x"{code[0x0000328b-0x00003288,1]}", -- 0x00003288
    x"{code[0x0000328f-0x0000328c,1]}", -- 0x0000328c
    x"{code[0x00003293-0x00003290,1]}", -- 0x00003290
    x"{code[0x00003297-0x00003294,1]}", -- 0x00003294
    x"{code[0x0000329b-0x00003298,1]}", -- 0x00003298
    x"{code[0x0000329f-0x0000329c,1]}", -- 0x0000329c
    x"{code[0x000032a3-0x000032a0,1]}", -- 0x000032a0
    x"{code[0x000032a7-0x000032a4,1]}", -- 0x000032a4
    x"{code[0x000032ab-0x000032a8,1]}", -- 0x000032a8
    x"{code[0x000032af-0x000032ac,1]}", -- 0x000032ac
    x"{code[0x000032b3-0x000032b0,1]}", -- 0x000032b0
    x"{code[0x000032b7-0x000032b4,1]}", -- 0x000032b4
    x"{code[0x000032bb-0x000032b8,1]}", -- 0x000032b8
    x"{code[0x000032bf-0x000032bc,1]}", -- 0x000032bc
    x"{code[0x000032c3-0x000032c0,1]}", -- 0x000032c0
    x"{code[0x000032c7-0x000032c4,1]}", -- 0x000032c4
    x"{code[0x000032cb-0x000032c8,1]}", -- 0x000032c8
    x"{code[0x000032cf-0x000032cc,1]}", -- 0x000032cc
    x"{code[0x000032d3-0x000032d0,1]}", -- 0x000032d0
    x"{code[0x000032d7-0x000032d4,1]}", -- 0x000032d4
    x"{code[0x000032db-0x000032d8,1]}", -- 0x000032d8
    x"{code[0x000032df-0x000032dc,1]}", -- 0x000032dc
    x"{code[0x000032e3-0x000032e0,1]}", -- 0x000032e0
    x"{code[0x000032e7-0x000032e4,1]}", -- 0x000032e4
    x"{code[0x000032eb-0x000032e8,1]}", -- 0x000032e8
    x"{code[0x000032ef-0x000032ec,1]}", -- 0x000032ec
    x"{code[0x000032f3-0x000032f0,1]}", -- 0x000032f0
    x"{code[0x000032f7-0x000032f4,1]}", -- 0x000032f4
    x"{code[0x000032fb-0x000032f8,1]}", -- 0x000032f8
    x"{code[0x000032ff-0x000032fc,1]}", -- 0x000032fc
    x"{code[0x00003303-0x00003300,1]}", -- 0x00003300
    x"{code[0x00003307-0x00003304,1]}", -- 0x00003304
    x"{code[0x0000330b-0x00003308,1]}", -- 0x00003308
    x"{code[0x0000330f-0x0000330c,1]}", -- 0x0000330c
    x"{code[0x00003313-0x00003310,1]}", -- 0x00003310
    x"{code[0x00003317-0x00003314,1]}", -- 0x00003314
    x"{code[0x0000331b-0x00003318,1]}", -- 0x00003318
    x"{code[0x0000331f-0x0000331c,1]}", -- 0x0000331c
    x"{code[0x00003323-0x00003320,1]}", -- 0x00003320
    x"{code[0x00003327-0x00003324,1]}", -- 0x00003324
    x"{code[0x0000332b-0x00003328,1]}", -- 0x00003328
    x"{code[0x0000332f-0x0000332c,1]}", -- 0x0000332c
    x"{code[0x00003333-0x00003330,1]}", -- 0x00003330
    x"{code[0x00003337-0x00003334,1]}", -- 0x00003334
    x"{code[0x0000333b-0x00003338,1]}", -- 0x00003338
    x"{code[0x0000333f-0x0000333c,1]}", -- 0x0000333c
    x"{code[0x00003343-0x00003340,1]}", -- 0x00003340
    x"{code[0x00003347-0x00003344,1]}", -- 0x00003344
    x"{code[0x0000334b-0x00003348,1]}", -- 0x00003348
    x"{code[0x0000334f-0x0000334c,1]}", -- 0x0000334c
    x"{code[0x00003353-0x00003350,1]}", -- 0x00003350
    x"{code[0x00003357-0x00003354,1]}", -- 0x00003354
    x"{code[0x0000335b-0x00003358,1]}", -- 0x00003358
    x"{code[0x0000335f-0x0000335c,1]}", -- 0x0000335c
    x"{code[0x00003363-0x00003360,1]}", -- 0x00003360
    x"{code[0x00003367-0x00003364,1]}", -- 0x00003364
    x"{code[0x0000336b-0x00003368,1]}", -- 0x00003368
    x"{code[0x0000336f-0x0000336c,1]}", -- 0x0000336c
    x"{code[0x00003373-0x00003370,1]}", -- 0x00003370
    x"{code[0x00003377-0x00003374,1]}", -- 0x00003374
    x"{code[0x0000337b-0x00003378,1]}", -- 0x00003378
    x"{code[0x0000337f-0x0000337c,1]}", -- 0x0000337c
    x"{code[0x00003383-0x00003380,1]}", -- 0x00003380
    x"{code[0x00003387-0x00003384,1]}", -- 0x00003384
    x"{code[0x0000338b-0x00003388,1]}", -- 0x00003388
    x"{code[0x0000338f-0x0000338c,1]}", -- 0x0000338c
    x"{code[0x00003393-0x00003390,1]}", -- 0x00003390
    x"{code[0x00003397-0x00003394,1]}", -- 0x00003394
    x"{code[0x0000339b-0x00003398,1]}", -- 0x00003398
    x"{code[0x0000339f-0x0000339c,1]}", -- 0x0000339c
    x"{code[0x000033a3-0x000033a0,1]}", -- 0x000033a0
    x"{code[0x000033a7-0x000033a4,1]}", -- 0x000033a4
    x"{code[0x000033ab-0x000033a8,1]}", -- 0x000033a8
    x"{code[0x000033af-0x000033ac,1]}", -- 0x000033ac
    x"{code[0x000033b3-0x000033b0,1]}", -- 0x000033b0
    x"{code[0x000033b7-0x000033b4,1]}", -- 0x000033b4
    x"{code[0x000033bb-0x000033b8,1]}", -- 0x000033b8
    x"{code[0x000033bf-0x000033bc,1]}", -- 0x000033bc
    x"{code[0x000033c3-0x000033c0,1]}", -- 0x000033c0
    x"{code[0x000033c7-0x000033c4,1]}", -- 0x000033c4
    x"{code[0x000033cb-0x000033c8,1]}", -- 0x000033c8
    x"{code[0x000033cf-0x000033cc,1]}", -- 0x000033cc
    x"{code[0x000033d3-0x000033d0,1]}", -- 0x000033d0
    x"{code[0x000033d7-0x000033d4,1]}", -- 0x000033d4
    x"{code[0x000033db-0x000033d8,1]}", -- 0x000033d8
    x"{code[0x000033df-0x000033dc,1]}", -- 0x000033dc
    x"{code[0x000033e3-0x000033e0,1]}", -- 0x000033e0
    x"{code[0x000033e7-0x000033e4,1]}", -- 0x000033e4
    x"{code[0x000033eb-0x000033e8,1]}", -- 0x000033e8
    x"{code[0x000033ef-0x000033ec,1]}", -- 0x000033ec
    x"{code[0x000033f3-0x000033f0,1]}", -- 0x000033f0
    x"{code[0x000033f7-0x000033f4,1]}", -- 0x000033f4
    x"{code[0x000033fb-0x000033f8,1]}", -- 0x000033f8
    x"{code[0x000033ff-0x000033fc,1]}", -- 0x000033fc
    x"{code[0x00003403-0x00003400,1]}", -- 0x00003400
    x"{code[0x00003407-0x00003404,1]}", -- 0x00003404
    x"{code[0x0000340b-0x00003408,1]}", -- 0x00003408
    x"{code[0x0000340f-0x0000340c,1]}", -- 0x0000340c
    x"{code[0x00003413-0x00003410,1]}", -- 0x00003410
    x"{code[0x00003417-0x00003414,1]}", -- 0x00003414
    x"{code[0x0000341b-0x00003418,1]}", -- 0x00003418
    x"{code[0x0000341f-0x0000341c,1]}", -- 0x0000341c
    x"{code[0x00003423-0x00003420,1]}", -- 0x00003420
    x"{code[0x00003427-0x00003424,1]}", -- 0x00003424
    x"{code[0x0000342b-0x00003428,1]}", -- 0x00003428
    x"{code[0x0000342f-0x0000342c,1]}", -- 0x0000342c
    x"{code[0x00003433-0x00003430,1]}", -- 0x00003430
    x"{code[0x00003437-0x00003434,1]}", -- 0x00003434
    x"{code[0x0000343b-0x00003438,1]}", -- 0x00003438
    x"{code[0x0000343f-0x0000343c,1]}", -- 0x0000343c
    x"{code[0x00003443-0x00003440,1]}", -- 0x00003440
    x"{code[0x00003447-0x00003444,1]}", -- 0x00003444
    x"{code[0x0000344b-0x00003448,1]}", -- 0x00003448
    x"{code[0x0000344f-0x0000344c,1]}", -- 0x0000344c
    x"{code[0x00003453-0x00003450,1]}", -- 0x00003450
    x"{code[0x00003457-0x00003454,1]}", -- 0x00003454
    x"{code[0x0000345b-0x00003458,1]}", -- 0x00003458
    x"{code[0x0000345f-0x0000345c,1]}", -- 0x0000345c
    x"{code[0x00003463-0x00003460,1]}", -- 0x00003460
    x"{code[0x00003467-0x00003464,1]}", -- 0x00003464
    x"{code[0x0000346b-0x00003468,1]}", -- 0x00003468
    x"{code[0x0000346f-0x0000346c,1]}", -- 0x0000346c
    x"{code[0x00003473-0x00003470,1]}", -- 0x00003470
    x"{code[0x00003477-0x00003474,1]}", -- 0x00003474
    x"{code[0x0000347b-0x00003478,1]}", -- 0x00003478
    x"{code[0x0000347f-0x0000347c,1]}", -- 0x0000347c
    x"{code[0x00003483-0x00003480,1]}", -- 0x00003480
    x"{code[0x00003487-0x00003484,1]}", -- 0x00003484
    x"{code[0x0000348b-0x00003488,1]}", -- 0x00003488
    x"{code[0x0000348f-0x0000348c,1]}", -- 0x0000348c
    x"{code[0x00003493-0x00003490,1]}", -- 0x00003490
    x"{code[0x00003497-0x00003494,1]}", -- 0x00003494
    x"{code[0x0000349b-0x00003498,1]}", -- 0x00003498
    x"{code[0x0000349f-0x0000349c,1]}", -- 0x0000349c
    x"{code[0x000034a3-0x000034a0,1]}", -- 0x000034a0
    x"{code[0x000034a7-0x000034a4,1]}", -- 0x000034a4
    x"{code[0x000034ab-0x000034a8,1]}", -- 0x000034a8
    x"{code[0x000034af-0x000034ac,1]}", -- 0x000034ac
    x"{code[0x000034b3-0x000034b0,1]}", -- 0x000034b0
    x"{code[0x000034b7-0x000034b4,1]}", -- 0x000034b4
    x"{code[0x000034bb-0x000034b8,1]}", -- 0x000034b8
    x"{code[0x000034bf-0x000034bc,1]}", -- 0x000034bc
    x"{code[0x000034c3-0x000034c0,1]}", -- 0x000034c0
    x"{code[0x000034c7-0x000034c4,1]}", -- 0x000034c4
    x"{code[0x000034cb-0x000034c8,1]}", -- 0x000034c8
    x"{code[0x000034cf-0x000034cc,1]}", -- 0x000034cc
    x"{code[0x000034d3-0x000034d0,1]}", -- 0x000034d0
    x"{code[0x000034d7-0x000034d4,1]}", -- 0x000034d4
    x"{code[0x000034db-0x000034d8,1]}", -- 0x000034d8
    x"{code[0x000034df-0x000034dc,1]}", -- 0x000034dc
    x"{code[0x000034e3-0x000034e0,1]}", -- 0x000034e0
    x"{code[0x000034e7-0x000034e4,1]}", -- 0x000034e4
    x"{code[0x000034eb-0x000034e8,1]}", -- 0x000034e8
    x"{code[0x000034ef-0x000034ec,1]}", -- 0x000034ec
    x"{code[0x000034f3-0x000034f0,1]}", -- 0x000034f0
    x"{code[0x000034f7-0x000034f4,1]}", -- 0x000034f4
    x"{code[0x000034fb-0x000034f8,1]}", -- 0x000034f8
    x"{code[0x000034ff-0x000034fc,1]}", -- 0x000034fc
    x"{code[0x00003503-0x00003500,1]}", -- 0x00003500
    x"{code[0x00003507-0x00003504,1]}", -- 0x00003504
    x"{code[0x0000350b-0x00003508,1]}", -- 0x00003508
    x"{code[0x0000350f-0x0000350c,1]}", -- 0x0000350c
    x"{code[0x00003513-0x00003510,1]}", -- 0x00003510
    x"{code[0x00003517-0x00003514,1]}", -- 0x00003514
    x"{code[0x0000351b-0x00003518,1]}", -- 0x00003518
    x"{code[0x0000351f-0x0000351c,1]}", -- 0x0000351c
    x"{code[0x00003523-0x00003520,1]}", -- 0x00003520
    x"{code[0x00003527-0x00003524,1]}", -- 0x00003524
    x"{code[0x0000352b-0x00003528,1]}", -- 0x00003528
    x"{code[0x0000352f-0x0000352c,1]}", -- 0x0000352c
    x"{code[0x00003533-0x00003530,1]}", -- 0x00003530
    x"{code[0x00003537-0x00003534,1]}", -- 0x00003534
    x"{code[0x0000353b-0x00003538,1]}", -- 0x00003538
    x"{code[0x0000353f-0x0000353c,1]}", -- 0x0000353c
    x"{code[0x00003543-0x00003540,1]}", -- 0x00003540
    x"{code[0x00003547-0x00003544,1]}", -- 0x00003544
    x"{code[0x0000354b-0x00003548,1]}", -- 0x00003548
    x"{code[0x0000354f-0x0000354c,1]}", -- 0x0000354c
    x"{code[0x00003553-0x00003550,1]}", -- 0x00003550
    x"{code[0x00003557-0x00003554,1]}", -- 0x00003554
    x"{code[0x0000355b-0x00003558,1]}", -- 0x00003558
    x"{code[0x0000355f-0x0000355c,1]}", -- 0x0000355c
    x"{code[0x00003563-0x00003560,1]}", -- 0x00003560
    x"{code[0x00003567-0x00003564,1]}", -- 0x00003564
    x"{code[0x0000356b-0x00003568,1]}", -- 0x00003568
    x"{code[0x0000356f-0x0000356c,1]}", -- 0x0000356c
    x"{code[0x00003573-0x00003570,1]}", -- 0x00003570
    x"{code[0x00003577-0x00003574,1]}", -- 0x00003574
    x"{code[0x0000357b-0x00003578,1]}", -- 0x00003578
    x"{code[0x0000357f-0x0000357c,1]}", -- 0x0000357c
    x"{code[0x00003583-0x00003580,1]}", -- 0x00003580
    x"{code[0x00003587-0x00003584,1]}", -- 0x00003584
    x"{code[0x0000358b-0x00003588,1]}", -- 0x00003588
    x"{code[0x0000358f-0x0000358c,1]}", -- 0x0000358c
    x"{code[0x00003593-0x00003590,1]}", -- 0x00003590
    x"{code[0x00003597-0x00003594,1]}", -- 0x00003594
    x"{code[0x0000359b-0x00003598,1]}", -- 0x00003598
    x"{code[0x0000359f-0x0000359c,1]}", -- 0x0000359c
    x"{code[0x000035a3-0x000035a0,1]}", -- 0x000035a0
    x"{code[0x000035a7-0x000035a4,1]}", -- 0x000035a4
    x"{code[0x000035ab-0x000035a8,1]}", -- 0x000035a8
    x"{code[0x000035af-0x000035ac,1]}", -- 0x000035ac
    x"{code[0x000035b3-0x000035b0,1]}", -- 0x000035b0
    x"{code[0x000035b7-0x000035b4,1]}", -- 0x000035b4
    x"{code[0x000035bb-0x000035b8,1]}", -- 0x000035b8
    x"{code[0x000035bf-0x000035bc,1]}", -- 0x000035bc
    x"{code[0x000035c3-0x000035c0,1]}", -- 0x000035c0
    x"{code[0x000035c7-0x000035c4,1]}", -- 0x000035c4
    x"{code[0x000035cb-0x000035c8,1]}", -- 0x000035c8
    x"{code[0x000035cf-0x000035cc,1]}", -- 0x000035cc
    x"{code[0x000035d3-0x000035d0,1]}", -- 0x000035d0
    x"{code[0x000035d7-0x000035d4,1]}", -- 0x000035d4
    x"{code[0x000035db-0x000035d8,1]}", -- 0x000035d8
    x"{code[0x000035df-0x000035dc,1]}", -- 0x000035dc
    x"{code[0x000035e3-0x000035e0,1]}", -- 0x000035e0
    x"{code[0x000035e7-0x000035e4,1]}", -- 0x000035e4
    x"{code[0x000035eb-0x000035e8,1]}", -- 0x000035e8
    x"{code[0x000035ef-0x000035ec,1]}", -- 0x000035ec
    x"{code[0x000035f3-0x000035f0,1]}", -- 0x000035f0
    x"{code[0x000035f7-0x000035f4,1]}", -- 0x000035f4
    x"{code[0x000035fb-0x000035f8,1]}", -- 0x000035f8
    x"{code[0x000035ff-0x000035fc,1]}", -- 0x000035fc
    x"{code[0x00003603-0x00003600,1]}", -- 0x00003600
    x"{code[0x00003607-0x00003604,1]}", -- 0x00003604
    x"{code[0x0000360b-0x00003608,1]}", -- 0x00003608
    x"{code[0x0000360f-0x0000360c,1]}", -- 0x0000360c
    x"{code[0x00003613-0x00003610,1]}", -- 0x00003610
    x"{code[0x00003617-0x00003614,1]}", -- 0x00003614
    x"{code[0x0000361b-0x00003618,1]}", -- 0x00003618
    x"{code[0x0000361f-0x0000361c,1]}", -- 0x0000361c
    x"{code[0x00003623-0x00003620,1]}", -- 0x00003620
    x"{code[0x00003627-0x00003624,1]}", -- 0x00003624
    x"{code[0x0000362b-0x00003628,1]}", -- 0x00003628
    x"{code[0x0000362f-0x0000362c,1]}", -- 0x0000362c
    x"{code[0x00003633-0x00003630,1]}", -- 0x00003630
    x"{code[0x00003637-0x00003634,1]}", -- 0x00003634
    x"{code[0x0000363b-0x00003638,1]}", -- 0x00003638
    x"{code[0x0000363f-0x0000363c,1]}", -- 0x0000363c
    x"{code[0x00003643-0x00003640,1]}", -- 0x00003640
    x"{code[0x00003647-0x00003644,1]}", -- 0x00003644
    x"{code[0x0000364b-0x00003648,1]}", -- 0x00003648
    x"{code[0x0000364f-0x0000364c,1]}", -- 0x0000364c
    x"{code[0x00003653-0x00003650,1]}", -- 0x00003650
    x"{code[0x00003657-0x00003654,1]}", -- 0x00003654
    x"{code[0x0000365b-0x00003658,1]}", -- 0x00003658
    x"{code[0x0000365f-0x0000365c,1]}", -- 0x0000365c
    x"{code[0x00003663-0x00003660,1]}", -- 0x00003660
    x"{code[0x00003667-0x00003664,1]}", -- 0x00003664
    x"{code[0x0000366b-0x00003668,1]}", -- 0x00003668
    x"{code[0x0000366f-0x0000366c,1]}", -- 0x0000366c
    x"{code[0x00003673-0x00003670,1]}", -- 0x00003670
    x"{code[0x00003677-0x00003674,1]}", -- 0x00003674
    x"{code[0x0000367b-0x00003678,1]}", -- 0x00003678
    x"{code[0x0000367f-0x0000367c,1]}", -- 0x0000367c
    x"{code[0x00003683-0x00003680,1]}", -- 0x00003680
    x"{code[0x00003687-0x00003684,1]}", -- 0x00003684
    x"{code[0x0000368b-0x00003688,1]}", -- 0x00003688
    x"{code[0x0000368f-0x0000368c,1]}", -- 0x0000368c
    x"{code[0x00003693-0x00003690,1]}", -- 0x00003690
    x"{code[0x00003697-0x00003694,1]}", -- 0x00003694
    x"{code[0x0000369b-0x00003698,1]}", -- 0x00003698
    x"{code[0x0000369f-0x0000369c,1]}", -- 0x0000369c
    x"{code[0x000036a3-0x000036a0,1]}", -- 0x000036a0
    x"{code[0x000036a7-0x000036a4,1]}", -- 0x000036a4
    x"{code[0x000036ab-0x000036a8,1]}", -- 0x000036a8
    x"{code[0x000036af-0x000036ac,1]}", -- 0x000036ac
    x"{code[0x000036b3-0x000036b0,1]}", -- 0x000036b0
    x"{code[0x000036b7-0x000036b4,1]}", -- 0x000036b4
    x"{code[0x000036bb-0x000036b8,1]}", -- 0x000036b8
    x"{code[0x000036bf-0x000036bc,1]}", -- 0x000036bc
    x"{code[0x000036c3-0x000036c0,1]}", -- 0x000036c0
    x"{code[0x000036c7-0x000036c4,1]}", -- 0x000036c4
    x"{code[0x000036cb-0x000036c8,1]}", -- 0x000036c8
    x"{code[0x000036cf-0x000036cc,1]}", -- 0x000036cc
    x"{code[0x000036d3-0x000036d0,1]}", -- 0x000036d0
    x"{code[0x000036d7-0x000036d4,1]}", -- 0x000036d4
    x"{code[0x000036db-0x000036d8,1]}", -- 0x000036d8
    x"{code[0x000036df-0x000036dc,1]}", -- 0x000036dc
    x"{code[0x000036e3-0x000036e0,1]}", -- 0x000036e0
    x"{code[0x000036e7-0x000036e4,1]}", -- 0x000036e4
    x"{code[0x000036eb-0x000036e8,1]}", -- 0x000036e8
    x"{code[0x000036ef-0x000036ec,1]}", -- 0x000036ec
    x"{code[0x000036f3-0x000036f0,1]}", -- 0x000036f0
    x"{code[0x000036f7-0x000036f4,1]}", -- 0x000036f4
    x"{code[0x000036fb-0x000036f8,1]}", -- 0x000036f8
    x"{code[0x000036ff-0x000036fc,1]}", -- 0x000036fc
    x"{code[0x00003703-0x00003700,1]}", -- 0x00003700
    x"{code[0x00003707-0x00003704,1]}", -- 0x00003704
    x"{code[0x0000370b-0x00003708,1]}", -- 0x00003708
    x"{code[0x0000370f-0x0000370c,1]}", -- 0x0000370c
    x"{code[0x00003713-0x00003710,1]}", -- 0x00003710
    x"{code[0x00003717-0x00003714,1]}", -- 0x00003714
    x"{code[0x0000371b-0x00003718,1]}", -- 0x00003718
    x"{code[0x0000371f-0x0000371c,1]}", -- 0x0000371c
    x"{code[0x00003723-0x00003720,1]}", -- 0x00003720
    x"{code[0x00003727-0x00003724,1]}", -- 0x00003724
    x"{code[0x0000372b-0x00003728,1]}", -- 0x00003728
    x"{code[0x0000372f-0x0000372c,1]}", -- 0x0000372c
    x"{code[0x00003733-0x00003730,1]}", -- 0x00003730
    x"{code[0x00003737-0x00003734,1]}", -- 0x00003734
    x"{code[0x0000373b-0x00003738,1]}", -- 0x00003738
    x"{code[0x0000373f-0x0000373c,1]}", -- 0x0000373c
    x"{code[0x00003743-0x00003740,1]}", -- 0x00003740
    x"{code[0x00003747-0x00003744,1]}", -- 0x00003744
    x"{code[0x0000374b-0x00003748,1]}", -- 0x00003748
    x"{code[0x0000374f-0x0000374c,1]}", -- 0x0000374c
    x"{code[0x00003753-0x00003750,1]}", -- 0x00003750
    x"{code[0x00003757-0x00003754,1]}", -- 0x00003754
    x"{code[0x0000375b-0x00003758,1]}", -- 0x00003758
    x"{code[0x0000375f-0x0000375c,1]}", -- 0x0000375c
    x"{code[0x00003763-0x00003760,1]}", -- 0x00003760
    x"{code[0x00003767-0x00003764,1]}", -- 0x00003764
    x"{code[0x0000376b-0x00003768,1]}", -- 0x00003768
    x"{code[0x0000376f-0x0000376c,1]}", -- 0x0000376c
    x"{code[0x00003773-0x00003770,1]}", -- 0x00003770
    x"{code[0x00003777-0x00003774,1]}", -- 0x00003774
    x"{code[0x0000377b-0x00003778,1]}", -- 0x00003778
    x"{code[0x0000377f-0x0000377c,1]}", -- 0x0000377c
    x"{code[0x00003783-0x00003780,1]}", -- 0x00003780
    x"{code[0x00003787-0x00003784,1]}", -- 0x00003784
    x"{code[0x0000378b-0x00003788,1]}", -- 0x00003788
    x"{code[0x0000378f-0x0000378c,1]}", -- 0x0000378c
    x"{code[0x00003793-0x00003790,1]}", -- 0x00003790
    x"{code[0x00003797-0x00003794,1]}", -- 0x00003794
    x"{code[0x0000379b-0x00003798,1]}", -- 0x00003798
    x"{code[0x0000379f-0x0000379c,1]}", -- 0x0000379c
    x"{code[0x000037a3-0x000037a0,1]}", -- 0x000037a0
    x"{code[0x000037a7-0x000037a4,1]}", -- 0x000037a4
    x"{code[0x000037ab-0x000037a8,1]}", -- 0x000037a8
    x"{code[0x000037af-0x000037ac,1]}", -- 0x000037ac
    x"{code[0x000037b3-0x000037b0,1]}", -- 0x000037b0
    x"{code[0x000037b7-0x000037b4,1]}", -- 0x000037b4
    x"{code[0x000037bb-0x000037b8,1]}", -- 0x000037b8
    x"{code[0x000037bf-0x000037bc,1]}", -- 0x000037bc
    x"{code[0x000037c3-0x000037c0,1]}", -- 0x000037c0
    x"{code[0x000037c7-0x000037c4,1]}", -- 0x000037c4
    x"{code[0x000037cb-0x000037c8,1]}", -- 0x000037c8
    x"{code[0x000037cf-0x000037cc,1]}", -- 0x000037cc
    x"{code[0x000037d3-0x000037d0,1]}", -- 0x000037d0
    x"{code[0x000037d7-0x000037d4,1]}", -- 0x000037d4
    x"{code[0x000037db-0x000037d8,1]}", -- 0x000037d8
    x"{code[0x000037df-0x000037dc,1]}", -- 0x000037dc
    x"{code[0x000037e3-0x000037e0,1]}", -- 0x000037e0
    x"{code[0x000037e7-0x000037e4,1]}", -- 0x000037e4
    x"{code[0x000037eb-0x000037e8,1]}", -- 0x000037e8
    x"{code[0x000037ef-0x000037ec,1]}", -- 0x000037ec
    x"{code[0x000037f3-0x000037f0,1]}", -- 0x000037f0
    x"{code[0x000037f7-0x000037f4,1]}", -- 0x000037f4
    x"{code[0x000037fb-0x000037f8,1]}", -- 0x000037f8
    x"{code[0x000037ff-0x000037fc,1]}", -- 0x000037fc
    x"{code[0x00003803-0x00003800,1]}", -- 0x00003800
    x"{code[0x00003807-0x00003804,1]}", -- 0x00003804
    x"{code[0x0000380b-0x00003808,1]}", -- 0x00003808
    x"{code[0x0000380f-0x0000380c,1]}", -- 0x0000380c
    x"{code[0x00003813-0x00003810,1]}", -- 0x00003810
    x"{code[0x00003817-0x00003814,1]}", -- 0x00003814
    x"{code[0x0000381b-0x00003818,1]}", -- 0x00003818
    x"{code[0x0000381f-0x0000381c,1]}", -- 0x0000381c
    x"{code[0x00003823-0x00003820,1]}", -- 0x00003820
    x"{code[0x00003827-0x00003824,1]}", -- 0x00003824
    x"{code[0x0000382b-0x00003828,1]}", -- 0x00003828
    x"{code[0x0000382f-0x0000382c,1]}", -- 0x0000382c
    x"{code[0x00003833-0x00003830,1]}", -- 0x00003830
    x"{code[0x00003837-0x00003834,1]}", -- 0x00003834
    x"{code[0x0000383b-0x00003838,1]}", -- 0x00003838
    x"{code[0x0000383f-0x0000383c,1]}", -- 0x0000383c
    x"{code[0x00003843-0x00003840,1]}", -- 0x00003840
    x"{code[0x00003847-0x00003844,1]}", -- 0x00003844
    x"{code[0x0000384b-0x00003848,1]}", -- 0x00003848
    x"{code[0x0000384f-0x0000384c,1]}", -- 0x0000384c
    x"{code[0x00003853-0x00003850,1]}", -- 0x00003850
    x"{code[0x00003857-0x00003854,1]}", -- 0x00003854
    x"{code[0x0000385b-0x00003858,1]}", -- 0x00003858
    x"{code[0x0000385f-0x0000385c,1]}", -- 0x0000385c
    x"{code[0x00003863-0x00003860,1]}", -- 0x00003860
    x"{code[0x00003867-0x00003864,1]}", -- 0x00003864
    x"{code[0x0000386b-0x00003868,1]}", -- 0x00003868
    x"{code[0x0000386f-0x0000386c,1]}", -- 0x0000386c
    x"{code[0x00003873-0x00003870,1]}", -- 0x00003870
    x"{code[0x00003877-0x00003874,1]}", -- 0x00003874
    x"{code[0x0000387b-0x00003878,1]}", -- 0x00003878
    x"{code[0x0000387f-0x0000387c,1]}", -- 0x0000387c
    x"{code[0x00003883-0x00003880,1]}", -- 0x00003880
    x"{code[0x00003887-0x00003884,1]}", -- 0x00003884
    x"{code[0x0000388b-0x00003888,1]}", -- 0x00003888
    x"{code[0x0000388f-0x0000388c,1]}", -- 0x0000388c
    x"{code[0x00003893-0x00003890,1]}", -- 0x00003890
    x"{code[0x00003897-0x00003894,1]}", -- 0x00003894
    x"{code[0x0000389b-0x00003898,1]}", -- 0x00003898
    x"{code[0x0000389f-0x0000389c,1]}", -- 0x0000389c
    x"{code[0x000038a3-0x000038a0,1]}", -- 0x000038a0
    x"{code[0x000038a7-0x000038a4,1]}", -- 0x000038a4
    x"{code[0x000038ab-0x000038a8,1]}", -- 0x000038a8
    x"{code[0x000038af-0x000038ac,1]}", -- 0x000038ac
    x"{code[0x000038b3-0x000038b0,1]}", -- 0x000038b0
    x"{code[0x000038b7-0x000038b4,1]}", -- 0x000038b4
    x"{code[0x000038bb-0x000038b8,1]}", -- 0x000038b8
    x"{code[0x000038bf-0x000038bc,1]}", -- 0x000038bc
    x"{code[0x000038c3-0x000038c0,1]}", -- 0x000038c0
    x"{code[0x000038c7-0x000038c4,1]}", -- 0x000038c4
    x"{code[0x000038cb-0x000038c8,1]}", -- 0x000038c8
    x"{code[0x000038cf-0x000038cc,1]}", -- 0x000038cc
    x"{code[0x000038d3-0x000038d0,1]}", -- 0x000038d0
    x"{code[0x000038d7-0x000038d4,1]}", -- 0x000038d4
    x"{code[0x000038db-0x000038d8,1]}", -- 0x000038d8
    x"{code[0x000038df-0x000038dc,1]}", -- 0x000038dc
    x"{code[0x000038e3-0x000038e0,1]}", -- 0x000038e0
    x"{code[0x000038e7-0x000038e4,1]}", -- 0x000038e4
    x"{code[0x000038eb-0x000038e8,1]}", -- 0x000038e8
    x"{code[0x000038ef-0x000038ec,1]}", -- 0x000038ec
    x"{code[0x000038f3-0x000038f0,1]}", -- 0x000038f0
    x"{code[0x000038f7-0x000038f4,1]}", -- 0x000038f4
    x"{code[0x000038fb-0x000038f8,1]}", -- 0x000038f8
    x"{code[0x000038ff-0x000038fc,1]}", -- 0x000038fc
    x"{code[0x00003903-0x00003900,1]}", -- 0x00003900
    x"{code[0x00003907-0x00003904,1]}", -- 0x00003904
    x"{code[0x0000390b-0x00003908,1]}", -- 0x00003908
    x"{code[0x0000390f-0x0000390c,1]}", -- 0x0000390c
    x"{code[0x00003913-0x00003910,1]}", -- 0x00003910
    x"{code[0x00003917-0x00003914,1]}", -- 0x00003914
    x"{code[0x0000391b-0x00003918,1]}", -- 0x00003918
    x"{code[0x0000391f-0x0000391c,1]}", -- 0x0000391c
    x"{code[0x00003923-0x00003920,1]}", -- 0x00003920
    x"{code[0x00003927-0x00003924,1]}", -- 0x00003924
    x"{code[0x0000392b-0x00003928,1]}", -- 0x00003928
    x"{code[0x0000392f-0x0000392c,1]}", -- 0x0000392c
    x"{code[0x00003933-0x00003930,1]}", -- 0x00003930
    x"{code[0x00003937-0x00003934,1]}", -- 0x00003934
    x"{code[0x0000393b-0x00003938,1]}", -- 0x00003938
    x"{code[0x0000393f-0x0000393c,1]}", -- 0x0000393c
    x"{code[0x00003943-0x00003940,1]}", -- 0x00003940
    x"{code[0x00003947-0x00003944,1]}", -- 0x00003944
    x"{code[0x0000394b-0x00003948,1]}", -- 0x00003948
    x"{code[0x0000394f-0x0000394c,1]}", -- 0x0000394c
    x"{code[0x00003953-0x00003950,1]}", -- 0x00003950
    x"{code[0x00003957-0x00003954,1]}", -- 0x00003954
    x"{code[0x0000395b-0x00003958,1]}", -- 0x00003958
    x"{code[0x0000395f-0x0000395c,1]}", -- 0x0000395c
    x"{code[0x00003963-0x00003960,1]}", -- 0x00003960
    x"{code[0x00003967-0x00003964,1]}", -- 0x00003964
    x"{code[0x0000396b-0x00003968,1]}", -- 0x00003968
    x"{code[0x0000396f-0x0000396c,1]}", -- 0x0000396c
    x"{code[0x00003973-0x00003970,1]}", -- 0x00003970
    x"{code[0x00003977-0x00003974,1]}", -- 0x00003974
    x"{code[0x0000397b-0x00003978,1]}", -- 0x00003978
    x"{code[0x0000397f-0x0000397c,1]}", -- 0x0000397c
    x"{code[0x00003983-0x00003980,1]}", -- 0x00003980
    x"{code[0x00003987-0x00003984,1]}", -- 0x00003984
    x"{code[0x0000398b-0x00003988,1]}", -- 0x00003988
    x"{code[0x0000398f-0x0000398c,1]}", -- 0x0000398c
    x"{code[0x00003993-0x00003990,1]}", -- 0x00003990
    x"{code[0x00003997-0x00003994,1]}", -- 0x00003994
    x"{code[0x0000399b-0x00003998,1]}", -- 0x00003998
    x"{code[0x0000399f-0x0000399c,1]}", -- 0x0000399c
    x"{code[0x000039a3-0x000039a0,1]}", -- 0x000039a0
    x"{code[0x000039a7-0x000039a4,1]}", -- 0x000039a4
    x"{code[0x000039ab-0x000039a8,1]}", -- 0x000039a8
    x"{code[0x000039af-0x000039ac,1]}", -- 0x000039ac
    x"{code[0x000039b3-0x000039b0,1]}", -- 0x000039b0
    x"{code[0x000039b7-0x000039b4,1]}", -- 0x000039b4
    x"{code[0x000039bb-0x000039b8,1]}", -- 0x000039b8
    x"{code[0x000039bf-0x000039bc,1]}", -- 0x000039bc
    x"{code[0x000039c3-0x000039c0,1]}", -- 0x000039c0
    x"{code[0x000039c7-0x000039c4,1]}", -- 0x000039c4
    x"{code[0x000039cb-0x000039c8,1]}", -- 0x000039c8
    x"{code[0x000039cf-0x000039cc,1]}", -- 0x000039cc
    x"{code[0x000039d3-0x000039d0,1]}", -- 0x000039d0
    x"{code[0x000039d7-0x000039d4,1]}", -- 0x000039d4
    x"{code[0x000039db-0x000039d8,1]}", -- 0x000039d8
    x"{code[0x000039df-0x000039dc,1]}", -- 0x000039dc
    x"{code[0x000039e3-0x000039e0,1]}", -- 0x000039e0
    x"{code[0x000039e7-0x000039e4,1]}", -- 0x000039e4
    x"{code[0x000039eb-0x000039e8,1]}", -- 0x000039e8
    x"{code[0x000039ef-0x000039ec,1]}", -- 0x000039ec
    x"{code[0x000039f3-0x000039f0,1]}", -- 0x000039f0
    x"{code[0x000039f7-0x000039f4,1]}", -- 0x000039f4
    x"{code[0x000039fb-0x000039f8,1]}", -- 0x000039f8
    x"{code[0x000039ff-0x000039fc,1]}", -- 0x000039fc
    x"{code[0x00003a03-0x00003a00,1]}", -- 0x00003a00
    x"{code[0x00003a07-0x00003a04,1]}", -- 0x00003a04
    x"{code[0x00003a0b-0x00003a08,1]}", -- 0x00003a08
    x"{code[0x00003a0f-0x00003a0c,1]}", -- 0x00003a0c
    x"{code[0x00003a13-0x00003a10,1]}", -- 0x00003a10
    x"{code[0x00003a17-0x00003a14,1]}", -- 0x00003a14
    x"{code[0x00003a1b-0x00003a18,1]}", -- 0x00003a18
    x"{code[0x00003a1f-0x00003a1c,1]}", -- 0x00003a1c
    x"{code[0x00003a23-0x00003a20,1]}", -- 0x00003a20
    x"{code[0x00003a27-0x00003a24,1]}", -- 0x00003a24
    x"{code[0x00003a2b-0x00003a28,1]}", -- 0x00003a28
    x"{code[0x00003a2f-0x00003a2c,1]}", -- 0x00003a2c
    x"{code[0x00003a33-0x00003a30,1]}", -- 0x00003a30
    x"{code[0x00003a37-0x00003a34,1]}", -- 0x00003a34
    x"{code[0x00003a3b-0x00003a38,1]}", -- 0x00003a38
    x"{code[0x00003a3f-0x00003a3c,1]}", -- 0x00003a3c
    x"{code[0x00003a43-0x00003a40,1]}", -- 0x00003a40
    x"{code[0x00003a47-0x00003a44,1]}", -- 0x00003a44
    x"{code[0x00003a4b-0x00003a48,1]}", -- 0x00003a48
    x"{code[0x00003a4f-0x00003a4c,1]}", -- 0x00003a4c
    x"{code[0x00003a53-0x00003a50,1]}", -- 0x00003a50
    x"{code[0x00003a57-0x00003a54,1]}", -- 0x00003a54
    x"{code[0x00003a5b-0x00003a58,1]}", -- 0x00003a58
    x"{code[0x00003a5f-0x00003a5c,1]}", -- 0x00003a5c
    x"{code[0x00003a63-0x00003a60,1]}", -- 0x00003a60
    x"{code[0x00003a67-0x00003a64,1]}", -- 0x00003a64
    x"{code[0x00003a6b-0x00003a68,1]}", -- 0x00003a68
    x"{code[0x00003a6f-0x00003a6c,1]}", -- 0x00003a6c
    x"{code[0x00003a73-0x00003a70,1]}", -- 0x00003a70
    x"{code[0x00003a77-0x00003a74,1]}", -- 0x00003a74
    x"{code[0x00003a7b-0x00003a78,1]}", -- 0x00003a78
    x"{code[0x00003a7f-0x00003a7c,1]}", -- 0x00003a7c
    x"{code[0x00003a83-0x00003a80,1]}", -- 0x00003a80
    x"{code[0x00003a87-0x00003a84,1]}", -- 0x00003a84
    x"{code[0x00003a8b-0x00003a88,1]}", -- 0x00003a88
    x"{code[0x00003a8f-0x00003a8c,1]}", -- 0x00003a8c
    x"{code[0x00003a93-0x00003a90,1]}", -- 0x00003a90
    x"{code[0x00003a97-0x00003a94,1]}", -- 0x00003a94
    x"{code[0x00003a9b-0x00003a98,1]}", -- 0x00003a98
    x"{code[0x00003a9f-0x00003a9c,1]}", -- 0x00003a9c
    x"{code[0x00003aa3-0x00003aa0,1]}", -- 0x00003aa0
    x"{code[0x00003aa7-0x00003aa4,1]}", -- 0x00003aa4
    x"{code[0x00003aab-0x00003aa8,1]}", -- 0x00003aa8
    x"{code[0x00003aaf-0x00003aac,1]}", -- 0x00003aac
    x"{code[0x00003ab3-0x00003ab0,1]}", -- 0x00003ab0
    x"{code[0x00003ab7-0x00003ab4,1]}", -- 0x00003ab4
    x"{code[0x00003abb-0x00003ab8,1]}", -- 0x00003ab8
    x"{code[0x00003abf-0x00003abc,1]}", -- 0x00003abc
    x"{code[0x00003ac3-0x00003ac0,1]}", -- 0x00003ac0
    x"{code[0x00003ac7-0x00003ac4,1]}", -- 0x00003ac4
    x"{code[0x00003acb-0x00003ac8,1]}", -- 0x00003ac8
    x"{code[0x00003acf-0x00003acc,1]}", -- 0x00003acc
    x"{code[0x00003ad3-0x00003ad0,1]}", -- 0x00003ad0
    x"{code[0x00003ad7-0x00003ad4,1]}", -- 0x00003ad4
    x"{code[0x00003adb-0x00003ad8,1]}", -- 0x00003ad8
    x"{code[0x00003adf-0x00003adc,1]}", -- 0x00003adc
    x"{code[0x00003ae3-0x00003ae0,1]}", -- 0x00003ae0
    x"{code[0x00003ae7-0x00003ae4,1]}", -- 0x00003ae4
    x"{code[0x00003aeb-0x00003ae8,1]}", -- 0x00003ae8
    x"{code[0x00003aef-0x00003aec,1]}", -- 0x00003aec
    x"{code[0x00003af3-0x00003af0,1]}", -- 0x00003af0
    x"{code[0x00003af7-0x00003af4,1]}", -- 0x00003af4
    x"{code[0x00003afb-0x00003af8,1]}", -- 0x00003af8
    x"{code[0x00003aff-0x00003afc,1]}", -- 0x00003afc
    x"{code[0x00003b03-0x00003b00,1]}", -- 0x00003b00
    x"{code[0x00003b07-0x00003b04,1]}", -- 0x00003b04
    x"{code[0x00003b0b-0x00003b08,1]}", -- 0x00003b08
    x"{code[0x00003b0f-0x00003b0c,1]}", -- 0x00003b0c
    x"{code[0x00003b13-0x00003b10,1]}", -- 0x00003b10
    x"{code[0x00003b17-0x00003b14,1]}", -- 0x00003b14
    x"{code[0x00003b1b-0x00003b18,1]}", -- 0x00003b18
    x"{code[0x00003b1f-0x00003b1c,1]}", -- 0x00003b1c
    x"{code[0x00003b23-0x00003b20,1]}", -- 0x00003b20
    x"{code[0x00003b27-0x00003b24,1]}", -- 0x00003b24
    x"{code[0x00003b2b-0x00003b28,1]}", -- 0x00003b28
    x"{code[0x00003b2f-0x00003b2c,1]}", -- 0x00003b2c
    x"{code[0x00003b33-0x00003b30,1]}", -- 0x00003b30
    x"{code[0x00003b37-0x00003b34,1]}", -- 0x00003b34
    x"{code[0x00003b3b-0x00003b38,1]}", -- 0x00003b38
    x"{code[0x00003b3f-0x00003b3c,1]}", -- 0x00003b3c
    x"{code[0x00003b43-0x00003b40,1]}", -- 0x00003b40
    x"{code[0x00003b47-0x00003b44,1]}", -- 0x00003b44
    x"{code[0x00003b4b-0x00003b48,1]}", -- 0x00003b48
    x"{code[0x00003b4f-0x00003b4c,1]}", -- 0x00003b4c
    x"{code[0x00003b53-0x00003b50,1]}", -- 0x00003b50
    x"{code[0x00003b57-0x00003b54,1]}", -- 0x00003b54
    x"{code[0x00003b5b-0x00003b58,1]}", -- 0x00003b58
    x"{code[0x00003b5f-0x00003b5c,1]}", -- 0x00003b5c
    x"{code[0x00003b63-0x00003b60,1]}", -- 0x00003b60
    x"{code[0x00003b67-0x00003b64,1]}", -- 0x00003b64
    x"{code[0x00003b6b-0x00003b68,1]}", -- 0x00003b68
    x"{code[0x00003b6f-0x00003b6c,1]}", -- 0x00003b6c
    x"{code[0x00003b73-0x00003b70,1]}", -- 0x00003b70
    x"{code[0x00003b77-0x00003b74,1]}", -- 0x00003b74
    x"{code[0x00003b7b-0x00003b78,1]}", -- 0x00003b78
    x"{code[0x00003b7f-0x00003b7c,1]}", -- 0x00003b7c
    x"{code[0x00003b83-0x00003b80,1]}", -- 0x00003b80
    x"{code[0x00003b87-0x00003b84,1]}", -- 0x00003b84
    x"{code[0x00003b8b-0x00003b88,1]}", -- 0x00003b88
    x"{code[0x00003b8f-0x00003b8c,1]}", -- 0x00003b8c
    x"{code[0x00003b93-0x00003b90,1]}", -- 0x00003b90
    x"{code[0x00003b97-0x00003b94,1]}", -- 0x00003b94
    x"{code[0x00003b9b-0x00003b98,1]}", -- 0x00003b98
    x"{code[0x00003b9f-0x00003b9c,1]}", -- 0x00003b9c
    x"{code[0x00003ba3-0x00003ba0,1]}", -- 0x00003ba0
    x"{code[0x00003ba7-0x00003ba4,1]}", -- 0x00003ba4
    x"{code[0x00003bab-0x00003ba8,1]}", -- 0x00003ba8
    x"{code[0x00003baf-0x00003bac,1]}", -- 0x00003bac
    x"{code[0x00003bb3-0x00003bb0,1]}", -- 0x00003bb0
    x"{code[0x00003bb7-0x00003bb4,1]}", -- 0x00003bb4
    x"{code[0x00003bbb-0x00003bb8,1]}", -- 0x00003bb8
    x"{code[0x00003bbf-0x00003bbc,1]}", -- 0x00003bbc
    x"{code[0x00003bc3-0x00003bc0,1]}", -- 0x00003bc0
    x"{code[0x00003bc7-0x00003bc4,1]}", -- 0x00003bc4
    x"{code[0x00003bcb-0x00003bc8,1]}", -- 0x00003bc8
    x"{code[0x00003bcf-0x00003bcc,1]}", -- 0x00003bcc
    x"{code[0x00003bd3-0x00003bd0,1]}", -- 0x00003bd0
    x"{code[0x00003bd7-0x00003bd4,1]}", -- 0x00003bd4
    x"{code[0x00003bdb-0x00003bd8,1]}", -- 0x00003bd8
    x"{code[0x00003bdf-0x00003bdc,1]}", -- 0x00003bdc
    x"{code[0x00003be3-0x00003be0,1]}", -- 0x00003be0
    x"{code[0x00003be7-0x00003be4,1]}", -- 0x00003be4
    x"{code[0x00003beb-0x00003be8,1]}", -- 0x00003be8
    x"{code[0x00003bef-0x00003bec,1]}", -- 0x00003bec
    x"{code[0x00003bf3-0x00003bf0,1]}", -- 0x00003bf0
    x"{code[0x00003bf7-0x00003bf4,1]}", -- 0x00003bf4
    x"{code[0x00003bfb-0x00003bf8,1]}", -- 0x00003bf8
    x"{code[0x00003bff-0x00003bfc,1]}", -- 0x00003bfc
    x"{code[0x00003c03-0x00003c00,1]}", -- 0x00003c00
    x"{code[0x00003c07-0x00003c04,1]}", -- 0x00003c04
    x"{code[0x00003c0b-0x00003c08,1]}", -- 0x00003c08
    x"{code[0x00003c0f-0x00003c0c,1]}", -- 0x00003c0c
    x"{code[0x00003c13-0x00003c10,1]}", -- 0x00003c10
    x"{code[0x00003c17-0x00003c14,1]}", -- 0x00003c14
    x"{code[0x00003c1b-0x00003c18,1]}", -- 0x00003c18
    x"{code[0x00003c1f-0x00003c1c,1]}", -- 0x00003c1c
    x"{code[0x00003c23-0x00003c20,1]}", -- 0x00003c20
    x"{code[0x00003c27-0x00003c24,1]}", -- 0x00003c24
    x"{code[0x00003c2b-0x00003c28,1]}", -- 0x00003c28
    x"{code[0x00003c2f-0x00003c2c,1]}", -- 0x00003c2c
    x"{code[0x00003c33-0x00003c30,1]}", -- 0x00003c30
    x"{code[0x00003c37-0x00003c34,1]}", -- 0x00003c34
    x"{code[0x00003c3b-0x00003c38,1]}", -- 0x00003c38
    x"{code[0x00003c3f-0x00003c3c,1]}", -- 0x00003c3c
    x"{code[0x00003c43-0x00003c40,1]}", -- 0x00003c40
    x"{code[0x00003c47-0x00003c44,1]}", -- 0x00003c44
    x"{code[0x00003c4b-0x00003c48,1]}", -- 0x00003c48
    x"{code[0x00003c4f-0x00003c4c,1]}", -- 0x00003c4c
    x"{code[0x00003c53-0x00003c50,1]}", -- 0x00003c50
    x"{code[0x00003c57-0x00003c54,1]}", -- 0x00003c54
    x"{code[0x00003c5b-0x00003c58,1]}", -- 0x00003c58
    x"{code[0x00003c5f-0x00003c5c,1]}", -- 0x00003c5c
    x"{code[0x00003c63-0x00003c60,1]}", -- 0x00003c60
    x"{code[0x00003c67-0x00003c64,1]}", -- 0x00003c64
    x"{code[0x00003c6b-0x00003c68,1]}", -- 0x00003c68
    x"{code[0x00003c6f-0x00003c6c,1]}", -- 0x00003c6c
    x"{code[0x00003c73-0x00003c70,1]}", -- 0x00003c70
    x"{code[0x00003c77-0x00003c74,1]}", -- 0x00003c74
    x"{code[0x00003c7b-0x00003c78,1]}", -- 0x00003c78
    x"{code[0x00003c7f-0x00003c7c,1]}", -- 0x00003c7c
    x"{code[0x00003c83-0x00003c80,1]}", -- 0x00003c80
    x"{code[0x00003c87-0x00003c84,1]}", -- 0x00003c84
    x"{code[0x00003c8b-0x00003c88,1]}", -- 0x00003c88
    x"{code[0x00003c8f-0x00003c8c,1]}", -- 0x00003c8c
    x"{code[0x00003c93-0x00003c90,1]}", -- 0x00003c90
    x"{code[0x00003c97-0x00003c94,1]}", -- 0x00003c94
    x"{code[0x00003c9b-0x00003c98,1]}", -- 0x00003c98
    x"{code[0x00003c9f-0x00003c9c,1]}", -- 0x00003c9c
    x"{code[0x00003ca3-0x00003ca0,1]}", -- 0x00003ca0
    x"{code[0x00003ca7-0x00003ca4,1]}", -- 0x00003ca4
    x"{code[0x00003cab-0x00003ca8,1]}", -- 0x00003ca8
    x"{code[0x00003caf-0x00003cac,1]}", -- 0x00003cac
    x"{code[0x00003cb3-0x00003cb0,1]}", -- 0x00003cb0
    x"{code[0x00003cb7-0x00003cb4,1]}", -- 0x00003cb4
    x"{code[0x00003cbb-0x00003cb8,1]}", -- 0x00003cb8
    x"{code[0x00003cbf-0x00003cbc,1]}", -- 0x00003cbc
    x"{code[0x00003cc3-0x00003cc0,1]}", -- 0x00003cc0
    x"{code[0x00003cc7-0x00003cc4,1]}", -- 0x00003cc4
    x"{code[0x00003ccb-0x00003cc8,1]}", -- 0x00003cc8
    x"{code[0x00003ccf-0x00003ccc,1]}", -- 0x00003ccc
    x"{code[0x00003cd3-0x00003cd0,1]}", -- 0x00003cd0
    x"{code[0x00003cd7-0x00003cd4,1]}", -- 0x00003cd4
    x"{code[0x00003cdb-0x00003cd8,1]}", -- 0x00003cd8
    x"{code[0x00003cdf-0x00003cdc,1]}", -- 0x00003cdc
    x"{code[0x00003ce3-0x00003ce0,1]}", -- 0x00003ce0
    x"{code[0x00003ce7-0x00003ce4,1]}", -- 0x00003ce4
    x"{code[0x00003ceb-0x00003ce8,1]}", -- 0x00003ce8
    x"{code[0x00003cef-0x00003cec,1]}", -- 0x00003cec
    x"{code[0x00003cf3-0x00003cf0,1]}", -- 0x00003cf0
    x"{code[0x00003cf7-0x00003cf4,1]}", -- 0x00003cf4
    x"{code[0x00003cfb-0x00003cf8,1]}", -- 0x00003cf8
    x"{code[0x00003cff-0x00003cfc,1]}", -- 0x00003cfc
    x"{code[0x00003d03-0x00003d00,1]}", -- 0x00003d00
    x"{code[0x00003d07-0x00003d04,1]}", -- 0x00003d04
    x"{code[0x00003d0b-0x00003d08,1]}", -- 0x00003d08
    x"{code[0x00003d0f-0x00003d0c,1]}", -- 0x00003d0c
    x"{code[0x00003d13-0x00003d10,1]}", -- 0x00003d10
    x"{code[0x00003d17-0x00003d14,1]}", -- 0x00003d14
    x"{code[0x00003d1b-0x00003d18,1]}", -- 0x00003d18
    x"{code[0x00003d1f-0x00003d1c,1]}", -- 0x00003d1c
    x"{code[0x00003d23-0x00003d20,1]}", -- 0x00003d20
    x"{code[0x00003d27-0x00003d24,1]}", -- 0x00003d24
    x"{code[0x00003d2b-0x00003d28,1]}", -- 0x00003d28
    x"{code[0x00003d2f-0x00003d2c,1]}", -- 0x00003d2c
    x"{code[0x00003d33-0x00003d30,1]}", -- 0x00003d30
    x"{code[0x00003d37-0x00003d34,1]}", -- 0x00003d34
    x"{code[0x00003d3b-0x00003d38,1]}", -- 0x00003d38
    x"{code[0x00003d3f-0x00003d3c,1]}", -- 0x00003d3c
    x"{code[0x00003d43-0x00003d40,1]}", -- 0x00003d40
    x"{code[0x00003d47-0x00003d44,1]}", -- 0x00003d44
    x"{code[0x00003d4b-0x00003d48,1]}", -- 0x00003d48
    x"{code[0x00003d4f-0x00003d4c,1]}", -- 0x00003d4c
    x"{code[0x00003d53-0x00003d50,1]}", -- 0x00003d50
    x"{code[0x00003d57-0x00003d54,1]}", -- 0x00003d54
    x"{code[0x00003d5b-0x00003d58,1]}", -- 0x00003d58
    x"{code[0x00003d5f-0x00003d5c,1]}", -- 0x00003d5c
    x"{code[0x00003d63-0x00003d60,1]}", -- 0x00003d60
    x"{code[0x00003d67-0x00003d64,1]}", -- 0x00003d64
    x"{code[0x00003d6b-0x00003d68,1]}", -- 0x00003d68
    x"{code[0x00003d6f-0x00003d6c,1]}", -- 0x00003d6c
    x"{code[0x00003d73-0x00003d70,1]}", -- 0x00003d70
    x"{code[0x00003d77-0x00003d74,1]}", -- 0x00003d74
    x"{code[0x00003d7b-0x00003d78,1]}", -- 0x00003d78
    x"{code[0x00003d7f-0x00003d7c,1]}", -- 0x00003d7c
    x"{code[0x00003d83-0x00003d80,1]}", -- 0x00003d80
    x"{code[0x00003d87-0x00003d84,1]}", -- 0x00003d84
    x"{code[0x00003d8b-0x00003d88,1]}", -- 0x00003d88
    x"{code[0x00003d8f-0x00003d8c,1]}", -- 0x00003d8c
    x"{code[0x00003d93-0x00003d90,1]}", -- 0x00003d90
    x"{code[0x00003d97-0x00003d94,1]}", -- 0x00003d94
    x"{code[0x00003d9b-0x00003d98,1]}", -- 0x00003d98
    x"{code[0x00003d9f-0x00003d9c,1]}", -- 0x00003d9c
    x"{code[0x00003da3-0x00003da0,1]}", -- 0x00003da0
    x"{code[0x00003da7-0x00003da4,1]}", -- 0x00003da4
    x"{code[0x00003dab-0x00003da8,1]}", -- 0x00003da8
    x"{code[0x00003daf-0x00003dac,1]}", -- 0x00003dac
    x"{code[0x00003db3-0x00003db0,1]}", -- 0x00003db0
    x"{code[0x00003db7-0x00003db4,1]}", -- 0x00003db4
    x"{code[0x00003dbb-0x00003db8,1]}", -- 0x00003db8
    x"{code[0x00003dbf-0x00003dbc,1]}", -- 0x00003dbc
    x"{code[0x00003dc3-0x00003dc0,1]}", -- 0x00003dc0
    x"{code[0x00003dc7-0x00003dc4,1]}", -- 0x00003dc4
    x"{code[0x00003dcb-0x00003dc8,1]}", -- 0x00003dc8
    x"{code[0x00003dcf-0x00003dcc,1]}", -- 0x00003dcc
    x"{code[0x00003dd3-0x00003dd0,1]}", -- 0x00003dd0
    x"{code[0x00003dd7-0x00003dd4,1]}", -- 0x00003dd4
    x"{code[0x00003ddb-0x00003dd8,1]}", -- 0x00003dd8
    x"{code[0x00003ddf-0x00003ddc,1]}", -- 0x00003ddc
    x"{code[0x00003de3-0x00003de0,1]}", -- 0x00003de0
    x"{code[0x00003de7-0x00003de4,1]}", -- 0x00003de4
    x"{code[0x00003deb-0x00003de8,1]}", -- 0x00003de8
    x"{code[0x00003def-0x00003dec,1]}", -- 0x00003dec
    x"{code[0x00003df3-0x00003df0,1]}", -- 0x00003df0
    x"{code[0x00003df7-0x00003df4,1]}", -- 0x00003df4
    x"{code[0x00003dfb-0x00003df8,1]}", -- 0x00003df8
    x"{code[0x00003dff-0x00003dfc,1]}", -- 0x00003dfc
    x"{code[0x00003e03-0x00003e00,1]}", -- 0x00003e00
    x"{code[0x00003e07-0x00003e04,1]}", -- 0x00003e04
    x"{code[0x00003e0b-0x00003e08,1]}", -- 0x00003e08
    x"{code[0x00003e0f-0x00003e0c,1]}", -- 0x00003e0c
    x"{code[0x00003e13-0x00003e10,1]}", -- 0x00003e10
    x"{code[0x00003e17-0x00003e14,1]}", -- 0x00003e14
    x"{code[0x00003e1b-0x00003e18,1]}", -- 0x00003e18
    x"{code[0x00003e1f-0x00003e1c,1]}", -- 0x00003e1c
    x"{code[0x00003e23-0x00003e20,1]}", -- 0x00003e20
    x"{code[0x00003e27-0x00003e24,1]}", -- 0x00003e24
    x"{code[0x00003e2b-0x00003e28,1]}", -- 0x00003e28
    x"{code[0x00003e2f-0x00003e2c,1]}", -- 0x00003e2c
    x"{code[0x00003e33-0x00003e30,1]}", -- 0x00003e30
    x"{code[0x00003e37-0x00003e34,1]}", -- 0x00003e34
    x"{code[0x00003e3b-0x00003e38,1]}", -- 0x00003e38
    x"{code[0x00003e3f-0x00003e3c,1]}", -- 0x00003e3c
    x"{code[0x00003e43-0x00003e40,1]}", -- 0x00003e40
    x"{code[0x00003e47-0x00003e44,1]}", -- 0x00003e44
    x"{code[0x00003e4b-0x00003e48,1]}", -- 0x00003e48
    x"{code[0x00003e4f-0x00003e4c,1]}", -- 0x00003e4c
    x"{code[0x00003e53-0x00003e50,1]}", -- 0x00003e50
    x"{code[0x00003e57-0x00003e54,1]}", -- 0x00003e54
    x"{code[0x00003e5b-0x00003e58,1]}", -- 0x00003e58
    x"{code[0x00003e5f-0x00003e5c,1]}", -- 0x00003e5c
    x"{code[0x00003e63-0x00003e60,1]}", -- 0x00003e60
    x"{code[0x00003e67-0x00003e64,1]}", -- 0x00003e64
    x"{code[0x00003e6b-0x00003e68,1]}", -- 0x00003e68
    x"{code[0x00003e6f-0x00003e6c,1]}", -- 0x00003e6c
    x"{code[0x00003e73-0x00003e70,1]}", -- 0x00003e70
    x"{code[0x00003e77-0x00003e74,1]}", -- 0x00003e74
    x"{code[0x00003e7b-0x00003e78,1]}", -- 0x00003e78
    x"{code[0x00003e7f-0x00003e7c,1]}", -- 0x00003e7c
    x"{code[0x00003e83-0x00003e80,1]}", -- 0x00003e80
    x"{code[0x00003e87-0x00003e84,1]}", -- 0x00003e84
    x"{code[0x00003e8b-0x00003e88,1]}", -- 0x00003e88
    x"{code[0x00003e8f-0x00003e8c,1]}", -- 0x00003e8c
    x"{code[0x00003e93-0x00003e90,1]}", -- 0x00003e90
    x"{code[0x00003e97-0x00003e94,1]}", -- 0x00003e94
    x"{code[0x00003e9b-0x00003e98,1]}", -- 0x00003e98
    x"{code[0x00003e9f-0x00003e9c,1]}", -- 0x00003e9c
    x"{code[0x00003ea3-0x00003ea0,1]}", -- 0x00003ea0
    x"{code[0x00003ea7-0x00003ea4,1]}", -- 0x00003ea4
    x"{code[0x00003eab-0x00003ea8,1]}", -- 0x00003ea8
    x"{code[0x00003eaf-0x00003eac,1]}", -- 0x00003eac
    x"{code[0x00003eb3-0x00003eb0,1]}", -- 0x00003eb0
    x"{code[0x00003eb7-0x00003eb4,1]}", -- 0x00003eb4
    x"{code[0x00003ebb-0x00003eb8,1]}", -- 0x00003eb8
    x"{code[0x00003ebf-0x00003ebc,1]}", -- 0x00003ebc
    x"{code[0x00003ec3-0x00003ec0,1]}", -- 0x00003ec0
    x"{code[0x00003ec7-0x00003ec4,1]}", -- 0x00003ec4
    x"{code[0x00003ecb-0x00003ec8,1]}", -- 0x00003ec8
    x"{code[0x00003ecf-0x00003ecc,1]}", -- 0x00003ecc
    x"{code[0x00003ed3-0x00003ed0,1]}", -- 0x00003ed0
    x"{code[0x00003ed7-0x00003ed4,1]}", -- 0x00003ed4
    x"{code[0x00003edb-0x00003ed8,1]}", -- 0x00003ed8
    x"{code[0x00003edf-0x00003edc,1]}", -- 0x00003edc
    x"{code[0x00003ee3-0x00003ee0,1]}", -- 0x00003ee0
    x"{code[0x00003ee7-0x00003ee4,1]}", -- 0x00003ee4
    x"{code[0x00003eeb-0x00003ee8,1]}", -- 0x00003ee8
    x"{code[0x00003eef-0x00003eec,1]}", -- 0x00003eec
    x"{code[0x00003ef3-0x00003ef0,1]}", -- 0x00003ef0
    x"{code[0x00003ef7-0x00003ef4,1]}", -- 0x00003ef4
    x"{code[0x00003efb-0x00003ef8,1]}", -- 0x00003ef8
    x"{code[0x00003eff-0x00003efc,1]}", -- 0x00003efc
    x"{code[0x00003f03-0x00003f00,1]}", -- 0x00003f00
    x"{code[0x00003f07-0x00003f04,1]}", -- 0x00003f04
    x"{code[0x00003f0b-0x00003f08,1]}", -- 0x00003f08
    x"{code[0x00003f0f-0x00003f0c,1]}", -- 0x00003f0c
    x"{code[0x00003f13-0x00003f10,1]}", -- 0x00003f10
    x"{code[0x00003f17-0x00003f14,1]}", -- 0x00003f14
    x"{code[0x00003f1b-0x00003f18,1]}", -- 0x00003f18
    x"{code[0x00003f1f-0x00003f1c,1]}", -- 0x00003f1c
    x"{code[0x00003f23-0x00003f20,1]}", -- 0x00003f20
    x"{code[0x00003f27-0x00003f24,1]}", -- 0x00003f24
    x"{code[0x00003f2b-0x00003f28,1]}", -- 0x00003f28
    x"{code[0x00003f2f-0x00003f2c,1]}", -- 0x00003f2c
    x"{code[0x00003f33-0x00003f30,1]}", -- 0x00003f30
    x"{code[0x00003f37-0x00003f34,1]}", -- 0x00003f34
    x"{code[0x00003f3b-0x00003f38,1]}", -- 0x00003f38
    x"{code[0x00003f3f-0x00003f3c,1]}", -- 0x00003f3c
    x"{code[0x00003f43-0x00003f40,1]}", -- 0x00003f40
    x"{code[0x00003f47-0x00003f44,1]}", -- 0x00003f44
    x"{code[0x00003f4b-0x00003f48,1]}", -- 0x00003f48
    x"{code[0x00003f4f-0x00003f4c,1]}", -- 0x00003f4c
    x"{code[0x00003f53-0x00003f50,1]}", -- 0x00003f50
    x"{code[0x00003f57-0x00003f54,1]}", -- 0x00003f54
    x"{code[0x00003f5b-0x00003f58,1]}", -- 0x00003f58
    x"{code[0x00003f5f-0x00003f5c,1]}", -- 0x00003f5c
    x"{code[0x00003f63-0x00003f60,1]}", -- 0x00003f60
    x"{code[0x00003f67-0x00003f64,1]}", -- 0x00003f64
    x"{code[0x00003f6b-0x00003f68,1]}", -- 0x00003f68
    x"{code[0x00003f6f-0x00003f6c,1]}", -- 0x00003f6c
    x"{code[0x00003f73-0x00003f70,1]}", -- 0x00003f70
    x"{code[0x00003f77-0x00003f74,1]}", -- 0x00003f74
    x"{code[0x00003f7b-0x00003f78,1]}", -- 0x00003f78
    x"{code[0x00003f7f-0x00003f7c,1]}", -- 0x00003f7c
    x"{code[0x00003f83-0x00003f80,1]}", -- 0x00003f80
    x"{code[0x00003f87-0x00003f84,1]}", -- 0x00003f84
    x"{code[0x00003f8b-0x00003f88,1]}", -- 0x00003f88
    x"{code[0x00003f8f-0x00003f8c,1]}", -- 0x00003f8c
    x"{code[0x00003f93-0x00003f90,1]}", -- 0x00003f90
    x"{code[0x00003f97-0x00003f94,1]}", -- 0x00003f94
    x"{code[0x00003f9b-0x00003f98,1]}", -- 0x00003f98
    x"{code[0x00003f9f-0x00003f9c,1]}", -- 0x00003f9c
    x"{code[0x00003fa3-0x00003fa0,1]}", -- 0x00003fa0
    x"{code[0x00003fa7-0x00003fa4,1]}", -- 0x00003fa4
    x"{code[0x00003fab-0x00003fa8,1]}", -- 0x00003fa8
    x"{code[0x00003faf-0x00003fac,1]}", -- 0x00003fac
    x"{code[0x00003fb3-0x00003fb0,1]}", -- 0x00003fb0
    x"{code[0x00003fb7-0x00003fb4,1]}", -- 0x00003fb4
    x"{code[0x00003fbb-0x00003fb8,1]}", -- 0x00003fb8
    x"{code[0x00003fbf-0x00003fbc,1]}", -- 0x00003fbc
    x"{code[0x00003fc3-0x00003fc0,1]}", -- 0x00003fc0
    x"{code[0x00003fc7-0x00003fc4,1]}", -- 0x00003fc4
    x"{code[0x00003fcb-0x00003fc8,1]}", -- 0x00003fc8
    x"{code[0x00003fcf-0x00003fcc,1]}", -- 0x00003fcc
    x"{code[0x00003fd3-0x00003fd0,1]}", -- 0x00003fd0
    x"{code[0x00003fd7-0x00003fd4,1]}", -- 0x00003fd4
    x"{code[0x00003fdb-0x00003fd8,1]}", -- 0x00003fd8
    x"{code[0x00003fdf-0x00003fdc,1]}", -- 0x00003fdc
    x"{code[0x00003fe3-0x00003fe0,1]}", -- 0x00003fe0
    x"{code[0x00003fe7-0x00003fe4,1]}", -- 0x00003fe4
    x"{code[0x00003feb-0x00003fe8,1]}", -- 0x00003fe8
    x"{code[0x00003fef-0x00003fec,1]}", -- 0x00003fec
    x"{code[0x00003ff3-0x00003ff0,1]}", -- 0x00003ff0
    x"{code[0x00003ff7-0x00003ff4,1]}", -- 0x00003ff4
    x"{code[0x00003ffb-0x00003ff8,1]}", -- 0x00003ff8
    x"{code[0x00003fff-0x00003ffc,1]}"  -- 0x00003ffc
  );
begin
  ACK_O <= read_ack or write_ack;
  DAT_O <= DAT_O_i;

  write_ack <= STB_I and WE_I;

  lookup_proc: process(CLK_I)
    variable addr : integer range 0 to 2 ** (ADR_I'length - 2) - 1;
  begin
    if rising_edge(CLK_I) then
      read_ack <= '0';
      DAT_O_i  <= (others=>'-');

      if RST_I = '0' then            
        if STB_I = '1' then 

          if WE_I = '0' and read_ack = '0' then
            addr  := to_integer(unsigned(ADR_I(ADR_I'length - 1 downto 2)));
            DAT_O_i  <= memory(addr);
            read_ack <= '1';
          elsif WE_I = '1' then
            addr  := to_integer(unsigned(ADR_I(ADR_I'length - 1 downto 2)));
            for i in 3 downto 0 loop
              if SEL_I(i) = '1' then
                memory(addr)(8 * i + 7 downto 8 * i) <= DAT_I(8 * i + 7 downto 8 * i);
              end if;
            end loop;
          end if;
        end if;
      end if;
    end if;
  end process;
end architecture;